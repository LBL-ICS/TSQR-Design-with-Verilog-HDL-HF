module multiplier(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [47:0] io_out_s
);
  assign io_out_s = io_in_a * io_in_b; // @[BinaryDesigns.scala 81:23]
endmodule
module full_subber(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s,
  output       io_out_c
);
  wire [8:0] _result_T = io_in_a - io_in_b; // @[BinaryDesigns.scala 69:23]
  wire [9:0] _result_T_2 = _result_T - 9'h0; // @[BinaryDesigns.scala 69:34]
  wire [8:0] result = _result_T_2[8:0]; // @[BinaryDesigns.scala 68:22 69:12]
  assign io_out_s = result[7:0]; // @[BinaryDesigns.scala 70:23]
  assign io_out_c = result[8]; // @[BinaryDesigns.scala 71:23]
endmodule
module twoscomplement(
  input  [7:0] io_in,
  output [7:0] io_out
);
  wire [7:0] _x_T = ~io_in; // @[BinaryDesigns.scala 25:16]
  assign io_out = 8'h1 + _x_T; // @[BinaryDesigns.scala 25:14]
endmodule
module full_adder(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s,
  output       io_out_c
);
  wire [8:0] _result_T = io_in_a + io_in_b; // @[BinaryDesigns.scala 55:23]
  wire [9:0] _result_T_1 = {{1'd0}, _result_T}; // @[BinaryDesigns.scala 55:34]
  wire [8:0] result = _result_T_1[8:0]; // @[BinaryDesigns.scala 54:22 55:12]
  assign io_out_s = result[7:0]; // @[BinaryDesigns.scala 56:23]
  assign io_out_c = result[8]; // @[BinaryDesigns.scala 57:23]
endmodule
module FP_multiplier_10ccs(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
`endif // RANDOMIZE_REG_INIT
  wire [23:0] multiplier_io_in_a; // @[FloatingPointDesigns.scala 1721:28]
  wire [23:0] multiplier_io_in_b; // @[FloatingPointDesigns.scala 1721:28]
  wire [47:0] multiplier_io_out_s; // @[FloatingPointDesigns.scala 1721:28]
  wire [7:0] subber_io_in_a; // @[FloatingPointDesigns.scala 1728:24]
  wire [7:0] subber_io_in_b; // @[FloatingPointDesigns.scala 1728:24]
  wire [7:0] subber_io_out_s; // @[FloatingPointDesigns.scala 1728:24]
  wire  subber_io_out_c; // @[FloatingPointDesigns.scala 1728:24]
  wire [7:0] complementN_io_in; // @[FloatingPointDesigns.scala 1737:29]
  wire [7:0] complementN_io_out; // @[FloatingPointDesigns.scala 1737:29]
  wire [7:0] adderN_io_in_a; // @[FloatingPointDesigns.scala 1754:24]
  wire [7:0] adderN_io_in_b; // @[FloatingPointDesigns.scala 1754:24]
  wire [7:0] adderN_io_out_s; // @[FloatingPointDesigns.scala 1754:24]
  wire  adderN_io_out_c; // @[FloatingPointDesigns.scala 1754:24]
  wire  s_0 = io_in_a[31]; // @[FloatingPointDesigns.scala 1687:20]
  wire  s_1 = io_in_b[31]; // @[FloatingPointDesigns.scala 1688:20]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FloatingPointDesigns.scala 1692:64]
  wire [8:0] _GEN_63 = {{1'd0}, io_in_a[30:23]}; // @[FloatingPointDesigns.scala 1692:36]
  wire [7:0] _GEN_0 = io_in_a[30:23] < 8'h1 ? 8'h1 : io_in_a[30:23]; // @[FloatingPointDesigns.scala 1694:45 1695:14 1697:14]
  wire [8:0] _GEN_1 = _GEN_63 > _T_2 ? _T_2 : {{1'd0}, _GEN_0}; // @[FloatingPointDesigns.scala 1692:71 1693:14]
  wire [8:0] _GEN_64 = {{1'd0}, io_in_b[30:23]}; // @[FloatingPointDesigns.scala 1699:36]
  wire [7:0] _GEN_2 = io_in_b[30:23] < 8'h1 ? 8'h1 : io_in_b[30:23]; // @[FloatingPointDesigns.scala 1701:45 1702:14 1704:14]
  wire [8:0] _GEN_3 = _GEN_64 > _T_2 ? _T_2 : {{1'd0}, _GEN_2}; // @[FloatingPointDesigns.scala 1699:71 1700:14]
  wire [22:0] frac_0 = io_in_a[22:0]; // @[FloatingPointDesigns.scala 1709:23]
  wire [22:0] frac_1 = io_in_b[22:0]; // @[FloatingPointDesigns.scala 1710:23]
  wire [23:0] new_frac_0 = {1'h1,frac_0}; // @[FloatingPointDesigns.scala 1714:24]
  wire [23:0] new_frac_1 = {1'h1,frac_1}; // @[FloatingPointDesigns.scala 1715:24]
  reg  s_reg_0_0; // @[FloatingPointDesigns.scala 1717:24]
  reg  s_reg_0_1; // @[FloatingPointDesigns.scala 1717:24]
  reg  s_reg_1_0; // @[FloatingPointDesigns.scala 1717:24]
  reg  s_reg_1_1; // @[FloatingPointDesigns.scala 1717:24]
  reg  s_reg_2_0; // @[FloatingPointDesigns.scala 1717:24]
  reg  s_reg_2_1; // @[FloatingPointDesigns.scala 1717:24]
  reg  s_reg_3_0; // @[FloatingPointDesigns.scala 1717:24]
  reg  s_reg_3_1; // @[FloatingPointDesigns.scala 1717:24]
  reg  s_reg_4_0; // @[FloatingPointDesigns.scala 1717:24]
  reg  s_reg_4_1; // @[FloatingPointDesigns.scala 1717:24]
  reg [7:0] exp_reg_0_0; // @[FloatingPointDesigns.scala 1718:26]
  reg [7:0] exp_reg_0_1; // @[FloatingPointDesigns.scala 1718:26]
  reg [7:0] exp_reg_1_0; // @[FloatingPointDesigns.scala 1718:26]
  reg [7:0] exp_reg_1_1; // @[FloatingPointDesigns.scala 1718:26]
  reg [7:0] exp_reg_2_0; // @[FloatingPointDesigns.scala 1718:26]
  reg [7:0] exp_reg_2_1; // @[FloatingPointDesigns.scala 1718:26]
  reg [7:0] exp_reg_3_0; // @[FloatingPointDesigns.scala 1718:26]
  reg [7:0] exp_reg_3_1; // @[FloatingPointDesigns.scala 1718:26]
  reg [7:0] exp_reg_4_0; // @[FloatingPointDesigns.scala 1718:26]
  reg [7:0] exp_reg_4_1; // @[FloatingPointDesigns.scala 1718:26]
  reg [7:0] exp_reg_5_0; // @[FloatingPointDesigns.scala 1718:26]
  reg [7:0] exp_reg_5_1; // @[FloatingPointDesigns.scala 1718:26]
  reg [7:0] exp_reg_6_0; // @[FloatingPointDesigns.scala 1718:26]
  reg [7:0] exp_reg_6_1; // @[FloatingPointDesigns.scala 1718:26]
  reg [7:0] exp_reg_7_0; // @[FloatingPointDesigns.scala 1718:26]
  reg [7:0] exp_reg_7_1; // @[FloatingPointDesigns.scala 1718:26]
  reg [7:0] exp_reg_8_0; // @[FloatingPointDesigns.scala 1718:26]
  reg [7:0] exp_reg_8_1; // @[FloatingPointDesigns.scala 1718:26]
  reg [23:0] new_frac_reg_0_0; // @[FloatingPointDesigns.scala 1719:31]
  reg [23:0] new_frac_reg_0_1; // @[FloatingPointDesigns.scala 1719:31]
  reg [23:0] new_frac_reg_1_0; // @[FloatingPointDesigns.scala 1719:31]
  reg [23:0] new_frac_reg_1_1; // @[FloatingPointDesigns.scala 1719:31]
  reg [47:0] multipplier_out_s_reg_0; // @[FloatingPointDesigns.scala 1725:40]
  reg [47:0] multipplier_out_s_reg_1; // @[FloatingPointDesigns.scala 1725:40]
  reg [47:0] multipplier_out_s_reg_2; // @[FloatingPointDesigns.scala 1725:40]
  reg [47:0] multipplier_out_s_reg_3; // @[FloatingPointDesigns.scala 1725:40]
  reg [47:0] multipplier_out_s_reg_4; // @[FloatingPointDesigns.scala 1725:40]
  reg [47:0] multipplier_out_s_reg_5; // @[FloatingPointDesigns.scala 1725:40]
  reg [7:0] subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1733:35]
  reg [7:0] complementN_out_reg_0; // @[FloatingPointDesigns.scala 1740:38]
  reg [7:0] complementN_out_reg_1; // @[FloatingPointDesigns.scala 1740:38]
  reg [7:0] complementN_out_reg_2; // @[FloatingPointDesigns.scala 1740:38]
  wire  new_s = s_reg_4_0 ^ s_reg_4_1; // @[FloatingPointDesigns.scala 1743:26]
  reg  new_s_reg_0; // @[FloatingPointDesigns.scala 1745:28]
  reg  new_s_reg_1; // @[FloatingPointDesigns.scala 1745:28]
  reg  new_s_reg_2; // @[FloatingPointDesigns.scala 1745:28]
  reg  new_s_reg_3; // @[FloatingPointDesigns.scala 1745:28]
  wire  is_exp1_neg_wire = exp_reg_5_1 < 8'h7f; // @[FloatingPointDesigns.scala 1748:40]
  reg  is_exp1_neg_reg_0; // @[FloatingPointDesigns.scala 1750:34]
  reg  is_exp1_neg_reg_1; // @[FloatingPointDesigns.scala 1750:34]
  wire [7:0] _adderN_io_in_a_T_1 = exp_reg_6_0 + 8'h1; // @[FloatingPointDesigns.scala 1758:39]
  reg [7:0] adderN_out_s_reg_0; // @[FloatingPointDesigns.scala 1765:35]
  reg  adderN_out_c_reg_0; // @[FloatingPointDesigns.scala 1766:35]
  reg [7:0] new_exp_reg_0; // @[FloatingPointDesigns.scala 1768:30]
  reg [22:0] new_mant_reg_0; // @[FloatingPointDesigns.scala 1769:31]
  reg [31:0] reg_out_s; // @[FloatingPointDesigns.scala 1771:28]
  wire  _new_exp_reg_0_T_1 = ~adderN_out_c_reg_0; // @[FloatingPointDesigns.scala 1775:55]
  wire [7:0] _new_exp_reg_0_T_2 = ~adderN_out_c_reg_0 ? 8'h1 : adderN_out_s_reg_0; // @[FloatingPointDesigns.scala 1775:54]
  wire  _new_exp_reg_0_T_5 = adderN_out_c_reg_0 | adderN_out_s_reg_0 > 8'hfe; // @[FloatingPointDesigns.scala 1775:142]
  wire [7:0] _new_exp_reg_0_T_6 = adderN_out_c_reg_0 | adderN_out_s_reg_0 > 8'hfe ? 8'hfe : adderN_out_s_reg_0; // @[FloatingPointDesigns.scala 1775:114]
  wire [7:0] _new_exp_reg_0_T_7 = is_exp1_neg_reg_1 ? _new_exp_reg_0_T_2 : _new_exp_reg_0_T_6; // @[FloatingPointDesigns.scala 1775:30]
  wire [31:0] _reg_out_s_T_1 = {new_s_reg_3,new_exp_reg_0,new_mant_reg_0}; // @[FloatingPointDesigns.scala 1817:53]
  wire [7:0] exp_0 = _GEN_1[7:0]; // @[FloatingPointDesigns.scala 1691:19]
  wire [7:0] exp_1 = _GEN_3[7:0]; // @[FloatingPointDesigns.scala 1691:19]
  wire [47:0] _GEN_17 = multiplier_io_out_s; // @[FloatingPointDesigns.scala 1773:19 1785:32 1725:40]
  wire [7:0] _GEN_18 = subber_io_out_s; // @[FloatingPointDesigns.scala 1773:19 1786:27 1733:35]
  wire [7:0] _GEN_20 = complementN_io_out; // @[FloatingPointDesigns.scala 1773:19 1788:30 1740:38]
  wire [7:0] _GEN_23 = adderN_io_out_s; // @[FloatingPointDesigns.scala 1773:19 1791:27 1765:35]
  wire  _GEN_24 = adderN_io_out_c; // @[FloatingPointDesigns.scala 1773:19 1792:27 1766:35]
  multiplier multiplier ( // @[FloatingPointDesigns.scala 1721:28]
    .io_in_a(multiplier_io_in_a),
    .io_in_b(multiplier_io_in_b),
    .io_out_s(multiplier_io_out_s)
  );
  full_subber subber ( // @[FloatingPointDesigns.scala 1728:24]
    .io_in_a(subber_io_in_a),
    .io_in_b(subber_io_in_b),
    .io_out_s(subber_io_out_s),
    .io_out_c(subber_io_out_c)
  );
  twoscomplement complementN ( // @[FloatingPointDesigns.scala 1737:29]
    .io_in(complementN_io_in),
    .io_out(complementN_io_out)
  );
  full_adder adderN ( // @[FloatingPointDesigns.scala 1754:24]
    .io_in_a(adderN_io_in_a),
    .io_in_b(adderN_io_in_b),
    .io_out_s(adderN_io_out_s),
    .io_out_c(adderN_io_out_c)
  );
  assign io_out_s = reg_out_s; // @[FloatingPointDesigns.scala 1820:14]
  assign multiplier_io_in_a = new_frac_reg_1_0; // @[FloatingPointDesigns.scala 1722:24]
  assign multiplier_io_in_b = new_frac_reg_1_1; // @[FloatingPointDesigns.scala 1723:24]
  assign subber_io_in_a = 8'h7f; // @[FloatingPointDesigns.scala 1729:20]
  assign subber_io_in_b = exp_reg_2_1; // @[FloatingPointDesigns.scala 1730:20]
  assign complementN_io_in = subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1738:23]
  assign adderN_io_in_a = multipplier_out_s_reg_4[47] ? _adderN_io_in_a_T_1 : exp_reg_6_0; // @[FloatingPointDesigns.scala 1757:70 1758:22 1761:22]
  assign adderN_io_in_b = complementN_out_reg_2; // @[FloatingPointDesigns.scala 1757:70 1759:22 1762:22]
  always @(posedge clock) begin
    if (reset) begin // @[FloatingPointDesigns.scala 1717:24]
      s_reg_0_0 <= 1'h0; // @[FloatingPointDesigns.scala 1717:24]
    end else begin
      s_reg_0_0 <= s_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1717:24]
      s_reg_0_1 <= 1'h0; // @[FloatingPointDesigns.scala 1717:24]
    end else begin
      s_reg_0_1 <= s_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1717:24]
      s_reg_1_0 <= 1'h0; // @[FloatingPointDesigns.scala 1717:24]
    end else begin
      s_reg_1_0 <= s_reg_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1717:24]
      s_reg_1_1 <= 1'h0; // @[FloatingPointDesigns.scala 1717:24]
    end else begin
      s_reg_1_1 <= s_reg_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1717:24]
      s_reg_2_0 <= 1'h0; // @[FloatingPointDesigns.scala 1717:24]
    end else begin
      s_reg_2_0 <= s_reg_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1717:24]
      s_reg_2_1 <= 1'h0; // @[FloatingPointDesigns.scala 1717:24]
    end else begin
      s_reg_2_1 <= s_reg_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1717:24]
      s_reg_3_0 <= 1'h0; // @[FloatingPointDesigns.scala 1717:24]
    end else begin
      s_reg_3_0 <= s_reg_2_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1717:24]
      s_reg_3_1 <= 1'h0; // @[FloatingPointDesigns.scala 1717:24]
    end else begin
      s_reg_3_1 <= s_reg_2_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1717:24]
      s_reg_4_0 <= 1'h0; // @[FloatingPointDesigns.scala 1717:24]
    end else begin
      s_reg_4_0 <= s_reg_3_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1717:24]
      s_reg_4_1 <= 1'h0; // @[FloatingPointDesigns.scala 1717:24]
    end else begin
      s_reg_4_1 <= s_reg_3_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_0_0 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_0_0 <= exp_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_0_1 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_0_1 <= exp_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_1_0 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_1_0 <= exp_reg_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_1_1 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_1_1 <= exp_reg_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_2_0 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_2_0 <= exp_reg_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_2_1 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_2_1 <= exp_reg_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_3_0 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_3_0 <= exp_reg_2_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_3_1 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_3_1 <= exp_reg_2_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_4_0 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_4_0 <= exp_reg_3_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_4_1 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_4_1 <= exp_reg_3_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_5_0 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_5_0 <= exp_reg_4_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_5_1 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_5_1 <= exp_reg_4_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_6_0 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_6_0 <= exp_reg_5_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_6_1 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_6_1 <= exp_reg_5_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_7_0 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_7_0 <= exp_reg_6_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_7_1 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_7_1 <= exp_reg_6_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_8_0 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_8_0 <= exp_reg_7_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1718:26]
      exp_reg_8_1 <= 8'h0; // @[FloatingPointDesigns.scala 1718:26]
    end else begin
      exp_reg_8_1 <= exp_reg_7_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1719:31]
      new_frac_reg_0_0 <= 24'h0; // @[FloatingPointDesigns.scala 1719:31]
    end else begin
      new_frac_reg_0_0 <= new_frac_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1719:31]
      new_frac_reg_0_1 <= 24'h0; // @[FloatingPointDesigns.scala 1719:31]
    end else begin
      new_frac_reg_0_1 <= new_frac_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1719:31]
      new_frac_reg_1_0 <= 24'h0; // @[FloatingPointDesigns.scala 1719:31]
    end else begin
      new_frac_reg_1_0 <= new_frac_reg_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1719:31]
      new_frac_reg_1_1 <= 24'h0; // @[FloatingPointDesigns.scala 1719:31]
    end else begin
      new_frac_reg_1_1 <= new_frac_reg_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1725:40]
      multipplier_out_s_reg_0 <= 48'h0; // @[FloatingPointDesigns.scala 1725:40]
    end else begin
      multipplier_out_s_reg_0 <= _GEN_17;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1725:40]
      multipplier_out_s_reg_1 <= 48'h0; // @[FloatingPointDesigns.scala 1725:40]
    end else begin
      multipplier_out_s_reg_1 <= multipplier_out_s_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1725:40]
      multipplier_out_s_reg_2 <= 48'h0; // @[FloatingPointDesigns.scala 1725:40]
    end else begin
      multipplier_out_s_reg_2 <= multipplier_out_s_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1725:40]
      multipplier_out_s_reg_3 <= 48'h0; // @[FloatingPointDesigns.scala 1725:40]
    end else begin
      multipplier_out_s_reg_3 <= multipplier_out_s_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1725:40]
      multipplier_out_s_reg_4 <= 48'h0; // @[FloatingPointDesigns.scala 1725:40]
    end else begin
      multipplier_out_s_reg_4 <= multipplier_out_s_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1725:40]
      multipplier_out_s_reg_5 <= 48'h0; // @[FloatingPointDesigns.scala 1725:40]
    end else begin
      multipplier_out_s_reg_5 <= multipplier_out_s_reg_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1733:35]
      subber_out_s_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1733:35]
    end else begin
      subber_out_s_reg_0 <= _GEN_18;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1740:38]
      complementN_out_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1740:38]
    end else begin
      complementN_out_reg_0 <= _GEN_20;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1740:38]
      complementN_out_reg_1 <= 8'h0; // @[FloatingPointDesigns.scala 1740:38]
    end else begin
      complementN_out_reg_1 <= complementN_out_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1740:38]
      complementN_out_reg_2 <= 8'h0; // @[FloatingPointDesigns.scala 1740:38]
    end else begin
      complementN_out_reg_2 <= complementN_out_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1745:28]
      new_s_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1745:28]
    end else begin
      new_s_reg_0 <= new_s;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1745:28]
      new_s_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1745:28]
    end else begin
      new_s_reg_1 <= new_s_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1745:28]
      new_s_reg_2 <= 1'h0; // @[FloatingPointDesigns.scala 1745:28]
    end else begin
      new_s_reg_2 <= new_s_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1745:28]
      new_s_reg_3 <= 1'h0; // @[FloatingPointDesigns.scala 1745:28]
    end else begin
      new_s_reg_3 <= new_s_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1750:34]
      is_exp1_neg_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1750:34]
    end else begin
      is_exp1_neg_reg_0 <= is_exp1_neg_wire;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1750:34]
      is_exp1_neg_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1750:34]
    end else begin
      is_exp1_neg_reg_1 <= is_exp1_neg_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1765:35]
      adderN_out_s_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1765:35]
    end else begin
      adderN_out_s_reg_0 <= _GEN_23;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1766:35]
      adderN_out_c_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1766:35]
    end else begin
      adderN_out_c_reg_0 <= _GEN_24;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1768:30]
      new_exp_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1768:30]
    end else if (multipplier_out_s_reg_5[47]) begin // @[FloatingPointDesigns.scala 1774:72]
      new_exp_reg_0 <= _new_exp_reg_0_T_7; // @[FloatingPointDesigns.scala 1775:24]
    end else begin
      new_exp_reg_0 <= _new_exp_reg_0_T_7; // @[FloatingPointDesigns.scala 1778:24]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1769:31]
      new_mant_reg_0 <= 23'h0; // @[FloatingPointDesigns.scala 1769:31]
    end else if (multipplier_out_s_reg_5[47]) begin // @[FloatingPointDesigns.scala 1774:72]
      if (is_exp1_neg_reg_1) begin // @[FloatingPointDesigns.scala 1776:31]
        if (_new_exp_reg_0_T_1) begin // @[FloatingPointDesigns.scala 1776:55]
          new_mant_reg_0 <= 23'h0;
        end else begin
          new_mant_reg_0 <= multipplier_out_s_reg_5[46:24];
        end
      end else if (_new_exp_reg_0_T_5) begin // @[FloatingPointDesigns.scala 1776:160]
        new_mant_reg_0 <= 23'h7fffff;
      end else begin
        new_mant_reg_0 <= multipplier_out_s_reg_5[46:24];
      end
    end else if (is_exp1_neg_reg_1) begin // @[FloatingPointDesigns.scala 1779:31]
      if (_new_exp_reg_0_T_1) begin // @[FloatingPointDesigns.scala 1779:55]
        new_mant_reg_0 <= 23'h0;
      end else begin
        new_mant_reg_0 <= multipplier_out_s_reg_5[45:23];
      end
    end else if (_new_exp_reg_0_T_5) begin // @[FloatingPointDesigns.scala 1779:156]
      new_mant_reg_0 <= 23'h7fffff;
    end else begin
      new_mant_reg_0 <= multipplier_out_s_reg_5[45:23];
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1771:28]
      reg_out_s <= 32'h0; // @[FloatingPointDesigns.scala 1771:28]
    end else if (exp_reg_8_0 == 8'h0 | exp_reg_8_1 == 8'h0) begin // @[FloatingPointDesigns.scala 1814:60]
      reg_out_s <= 32'h0; // @[FloatingPointDesigns.scala 1815:19]
    end else begin
      reg_out_s <= _reg_out_s_T_1; // @[FloatingPointDesigns.scala 1817:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s_reg_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s_reg_0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  s_reg_1_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  s_reg_1_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  s_reg_2_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  s_reg_2_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  s_reg_3_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  s_reg_3_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  s_reg_4_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  s_reg_4_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  exp_reg_0_0 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  exp_reg_0_1 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  exp_reg_1_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  exp_reg_1_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  exp_reg_2_0 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  exp_reg_2_1 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  exp_reg_3_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  exp_reg_3_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  exp_reg_4_0 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  exp_reg_4_1 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  exp_reg_5_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  exp_reg_5_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  exp_reg_6_0 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  exp_reg_6_1 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  exp_reg_7_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  exp_reg_7_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  exp_reg_8_0 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  exp_reg_8_1 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  new_frac_reg_0_0 = _RAND_28[23:0];
  _RAND_29 = {1{`RANDOM}};
  new_frac_reg_0_1 = _RAND_29[23:0];
  _RAND_30 = {1{`RANDOM}};
  new_frac_reg_1_0 = _RAND_30[23:0];
  _RAND_31 = {1{`RANDOM}};
  new_frac_reg_1_1 = _RAND_31[23:0];
  _RAND_32 = {2{`RANDOM}};
  multipplier_out_s_reg_0 = _RAND_32[47:0];
  _RAND_33 = {2{`RANDOM}};
  multipplier_out_s_reg_1 = _RAND_33[47:0];
  _RAND_34 = {2{`RANDOM}};
  multipplier_out_s_reg_2 = _RAND_34[47:0];
  _RAND_35 = {2{`RANDOM}};
  multipplier_out_s_reg_3 = _RAND_35[47:0];
  _RAND_36 = {2{`RANDOM}};
  multipplier_out_s_reg_4 = _RAND_36[47:0];
  _RAND_37 = {2{`RANDOM}};
  multipplier_out_s_reg_5 = _RAND_37[47:0];
  _RAND_38 = {1{`RANDOM}};
  subber_out_s_reg_0 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  complementN_out_reg_0 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  complementN_out_reg_1 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  complementN_out_reg_2 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  new_s_reg_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  new_s_reg_1 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  new_s_reg_2 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  new_s_reg_3 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  is_exp1_neg_reg_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  is_exp1_neg_reg_1 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  adderN_out_s_reg_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  adderN_out_c_reg_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  new_exp_reg_0 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  new_mant_reg_0 = _RAND_51[22:0];
  _RAND_52 = {1{`RANDOM}};
  reg_out_s = _RAND_52[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module full_adder_128(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [23:0] io_out_s,
  output        io_out_c
);
  wire [24:0] _result_T = io_in_a + io_in_b; // @[BinaryDesigns.scala 55:23]
  wire [25:0] _result_T_1 = {{1'd0}, _result_T}; // @[BinaryDesigns.scala 55:34]
  wire [24:0] result = _result_T_1[24:0]; // @[BinaryDesigns.scala 54:22 55:12]
  assign io_out_s = result[23:0]; // @[BinaryDesigns.scala 56:23]
  assign io_out_c = result[24]; // @[BinaryDesigns.scala 57:23]
endmodule
module FP_adder_13ccs(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] subber_io_in_a; // @[FloatingPointDesigns.scala 1456:24]
  wire [7:0] subber_io_in_b; // @[FloatingPointDesigns.scala 1456:24]
  wire [7:0] subber_io_out_s; // @[FloatingPointDesigns.scala 1456:24]
  wire  subber_io_out_c; // @[FloatingPointDesigns.scala 1456:24]
  wire [23:0] adder_io_in_a; // @[FloatingPointDesigns.scala 1462:23]
  wire [23:0] adder_io_in_b; // @[FloatingPointDesigns.scala 1462:23]
  wire [23:0] adder_io_out_s; // @[FloatingPointDesigns.scala 1462:23]
  wire  adder_io_out_c; // @[FloatingPointDesigns.scala 1462:23]
  wire [7:0] subber2_io_in_a; // @[FloatingPointDesigns.scala 1523:25]
  wire [7:0] subber2_io_in_b; // @[FloatingPointDesigns.scala 1523:25]
  wire [7:0] subber2_io_out_s; // @[FloatingPointDesigns.scala 1523:25]
  wire  subber2_io_out_c; // @[FloatingPointDesigns.scala 1523:25]
  wire  sign_0 = io_in_a[31]; // @[FloatingPointDesigns.scala 1385:23]
  wire  sign_1 = io_in_b[31]; // @[FloatingPointDesigns.scala 1386:23]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FloatingPointDesigns.scala 1389:64]
  wire [8:0] _GEN_167 = {{1'd0}, io_in_a[30:23]}; // @[FloatingPointDesigns.scala 1389:36]
  wire [7:0] _GEN_0 = io_in_a[30:23] < 8'h1 ? 8'h1 : io_in_a[30:23]; // @[FloatingPointDesigns.scala 1391:46 1392:14 1394:14]
  wire [8:0] _GEN_1 = _GEN_167 > _T_2 ? _T_2 : {{1'd0}, _GEN_0}; // @[FloatingPointDesigns.scala 1389:71 1390:14]
  wire [8:0] _GEN_168 = {{1'd0}, io_in_b[30:23]}; // @[FloatingPointDesigns.scala 1396:36]
  wire [7:0] _GEN_2 = io_in_b[30:23] < 8'h1 ? 8'h1 : io_in_b[30:23]; // @[FloatingPointDesigns.scala 1398:45 1399:14 1401:14]
  wire [8:0] _GEN_3 = _GEN_168 > _T_2 ? _T_2 : {{1'd0}, _GEN_2}; // @[FloatingPointDesigns.scala 1396:71 1397:14]
  wire [22:0] frac_0 = io_in_a[22:0]; // @[FloatingPointDesigns.scala 1406:23]
  wire [22:0] frac_1 = io_in_b[22:0]; // @[FloatingPointDesigns.scala 1407:23]
  wire [23:0] whole_frac_0 = {1'h1,frac_0}; // @[FloatingPointDesigns.scala 1411:26]
  wire [23:0] whole_frac_1 = {1'h1,frac_1}; // @[FloatingPointDesigns.scala 1412:26]
  reg  sign_reg_0_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_0_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_1_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_1_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_2_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_2_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_3_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_3_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_4_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_4_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_5_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_5_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_6_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_6_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_7_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_7_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_8_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_8_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_9_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_9_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_10_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_10_1; // @[FloatingPointDesigns.scala 1414:28]
  reg [7:0] exp_reg_0_0; // @[FloatingPointDesigns.scala 1415:28]
  reg [7:0] exp_reg_0_1; // @[FloatingPointDesigns.scala 1415:28]
  reg [7:0] exp_reg_1_0; // @[FloatingPointDesigns.scala 1415:28]
  reg [7:0] exp_reg_1_1; // @[FloatingPointDesigns.scala 1415:28]
  reg [7:0] exp_reg_2_0; // @[FloatingPointDesigns.scala 1415:28]
  reg [7:0] exp_reg_2_1; // @[FloatingPointDesigns.scala 1415:28]
  reg [22:0] frac_reg_0_0; // @[FloatingPointDesigns.scala 1416:28]
  reg [22:0] frac_reg_0_1; // @[FloatingPointDesigns.scala 1416:28]
  reg [22:0] frac_reg_1_0; // @[FloatingPointDesigns.scala 1416:28]
  reg [22:0] frac_reg_1_1; // @[FloatingPointDesigns.scala 1416:28]
  reg [22:0] frac_reg_2_0; // @[FloatingPointDesigns.scala 1416:28]
  reg [22:0] frac_reg_2_1; // @[FloatingPointDesigns.scala 1416:28]
  reg [23:0] wfrac_reg_0_0; // @[FloatingPointDesigns.scala 1417:28]
  reg [23:0] wfrac_reg_0_1; // @[FloatingPointDesigns.scala 1417:28]
  reg [23:0] wfrac_reg_1_0; // @[FloatingPointDesigns.scala 1417:28]
  reg [23:0] wfrac_reg_1_1; // @[FloatingPointDesigns.scala 1417:28]
  reg [23:0] wfrac_reg_2_0; // @[FloatingPointDesigns.scala 1417:28]
  reg [23:0] wfrac_reg_2_1; // @[FloatingPointDesigns.scala 1417:28]
  reg [7:0] subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1419:35]
  reg [7:0] subber_out_s_reg_1; // @[FloatingPointDesigns.scala 1419:35]
  reg  subber_out_c_reg_0; // @[FloatingPointDesigns.scala 1420:35]
  reg  subber_out_c_reg_1; // @[FloatingPointDesigns.scala 1420:35]
  reg [23:0] wire_temp_add_in_reg_0_0; // @[FloatingPointDesigns.scala 1422:39]
  reg [23:0] wire_temp_add_in_reg_0_1; // @[FloatingPointDesigns.scala 1422:39]
  reg [23:0] wire_temp_add_in_reg_1_0; // @[FloatingPointDesigns.scala 1422:39]
  reg [23:0] wire_temp_add_in_reg_1_1; // @[FloatingPointDesigns.scala 1422:39]
  reg  ref_s_reg_0; // @[FloatingPointDesigns.scala 1424:31]
  reg  ref_s_reg_1; // @[FloatingPointDesigns.scala 1424:31]
  reg  ref_s_reg_2; // @[FloatingPointDesigns.scala 1424:31]
  reg  ref_s_reg_3; // @[FloatingPointDesigns.scala 1424:31]
  reg  ref_s_reg_4; // @[FloatingPointDesigns.scala 1424:31]
  reg  ref_s_reg_5; // @[FloatingPointDesigns.scala 1424:31]
  reg  ref_s_reg_6; // @[FloatingPointDesigns.scala 1424:31]
  reg  ref_s_reg_7; // @[FloatingPointDesigns.scala 1424:31]
  reg [22:0] ref_frac_reg_0; // @[FloatingPointDesigns.scala 1425:31]
  reg [22:0] ref_frac_reg_1; // @[FloatingPointDesigns.scala 1425:31]
  reg [22:0] ref_frac_reg_2; // @[FloatingPointDesigns.scala 1425:31]
  reg [22:0] ref_frac_reg_3; // @[FloatingPointDesigns.scala 1425:31]
  reg [22:0] ref_frac_reg_4; // @[FloatingPointDesigns.scala 1425:31]
  reg [22:0] ref_frac_reg_5; // @[FloatingPointDesigns.scala 1425:31]
  reg [22:0] ref_frac_reg_6; // @[FloatingPointDesigns.scala 1425:31]
  reg [22:0] ref_frac_reg_7; // @[FloatingPointDesigns.scala 1425:31]
  reg [7:0] ref_exp_reg_0; // @[FloatingPointDesigns.scala 1426:31]
  reg [7:0] ref_exp_reg_1; // @[FloatingPointDesigns.scala 1426:31]
  reg [7:0] ref_exp_reg_2; // @[FloatingPointDesigns.scala 1426:31]
  reg [7:0] ref_exp_reg_3; // @[FloatingPointDesigns.scala 1426:31]
  reg [7:0] ref_exp_reg_4; // @[FloatingPointDesigns.scala 1426:31]
  reg [7:0] ref_exp_reg_5; // @[FloatingPointDesigns.scala 1426:31]
  reg [7:0] ref_exp_reg_6; // @[FloatingPointDesigns.scala 1426:31]
  reg [7:0] ref_exp_reg_7; // @[FloatingPointDesigns.scala 1426:31]
  reg [7:0] sub_exp_reg_0; // @[FloatingPointDesigns.scala 1427:31]
  reg [7:0] sub_exp_reg_1; // @[FloatingPointDesigns.scala 1427:31]
  reg [7:0] sub_exp_reg_2; // @[FloatingPointDesigns.scala 1427:31]
  reg [7:0] sub_exp_reg_3; // @[FloatingPointDesigns.scala 1427:31]
  reg [7:0] sub_exp_reg_4; // @[FloatingPointDesigns.scala 1427:31]
  reg [7:0] sub_exp_reg_5; // @[FloatingPointDesigns.scala 1427:31]
  reg [7:0] sub_exp_reg_6; // @[FloatingPointDesigns.scala 1427:31]
  reg [7:0] sub_exp_reg_7; // @[FloatingPointDesigns.scala 1427:31]
  reg [23:0] adder_io_out_s_reg_0; // @[FloatingPointDesigns.scala 1429:37]
  reg [23:0] adder_io_out_s_reg_1; // @[FloatingPointDesigns.scala 1429:37]
  reg [23:0] adder_io_out_s_reg_2; // @[FloatingPointDesigns.scala 1429:37]
  reg  adder_io_out_c_reg_0; // @[FloatingPointDesigns.scala 1430:37]
  reg  new_s_reg_0; // @[FloatingPointDesigns.scala 1432:35]
  reg  new_s_reg_1; // @[FloatingPointDesigns.scala 1432:35]
  reg  new_s_reg_2; // @[FloatingPointDesigns.scala 1432:35]
  reg  new_s_reg_3; // @[FloatingPointDesigns.scala 1432:35]
  reg  new_s_reg_4; // @[FloatingPointDesigns.scala 1432:35]
  reg  new_s_reg_5; // @[FloatingPointDesigns.scala 1432:35]
  reg [22:0] new_out_frac_reg_0; // @[FloatingPointDesigns.scala 1433:35]
  reg [7:0] new_out_exp_reg_0; // @[FloatingPointDesigns.scala 1434:35]
  reg  E_reg_0; // @[FloatingPointDesigns.scala 1435:24]
  reg  E_reg_1; // @[FloatingPointDesigns.scala 1435:24]
  reg  E_reg_2; // @[FloatingPointDesigns.scala 1435:24]
  reg  E_reg_3; // @[FloatingPointDesigns.scala 1435:24]
  reg  E_reg_4; // @[FloatingPointDesigns.scala 1435:24]
  reg  D_reg_0; // @[FloatingPointDesigns.scala 1436:24]
  reg  D_reg_1; // @[FloatingPointDesigns.scala 1436:24]
  reg  D_reg_2; // @[FloatingPointDesigns.scala 1436:24]
  reg  D_reg_3; // @[FloatingPointDesigns.scala 1436:24]
  reg  D_reg_4; // @[FloatingPointDesigns.scala 1436:24]
  reg [23:0] adder_result_reg_0; // @[FloatingPointDesigns.scala 1438:35]
  reg [23:0] adder_result_reg_1; // @[FloatingPointDesigns.scala 1438:35]
  reg [23:0] adder_result_reg_2; // @[FloatingPointDesigns.scala 1438:35]
  reg [5:0] leadingOne_reg_0; // @[FloatingPointDesigns.scala 1440:33]
  reg [5:0] leadingOne_reg_1; // @[FloatingPointDesigns.scala 1440:33]
  reg [31:0] io_in_a_reg_0; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_1; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_2; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_3; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_4; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_5; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_6; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_7; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_8; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_9; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_10; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_b_reg_0; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_1; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_2; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_3; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_4; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_5; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_6; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_7; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_8; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_9; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_10; // @[FloatingPointDesigns.scala 1443:30]
  reg [7:0] subber2_out_s_reg_0; // @[FloatingPointDesigns.scala 1445:36]
  reg  subber2_out_c_reg_0; // @[FloatingPointDesigns.scala 1446:36]
  reg [7:0] cmpl_subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1467:40]
  wire [7:0] _cmpl_subber_out_s_reg_0_T = ~subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1469:41]
  wire [7:0] _cmpl_subber_out_s_reg_0_T_2 = 8'h1 + _cmpl_subber_out_s_reg_0_T; // @[FloatingPointDesigns.scala 1469:39]
  wire [23:0] _wire_temp_add_in_0_T = wfrac_reg_2_0 >> cmpl_subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1477:46]
  wire [23:0] _wire_temp_add_in_1_T = wfrac_reg_2_1 >> subber_out_s_reg_1; // @[FloatingPointDesigns.scala 1485:46]
  reg [23:0] cmpl_wire_temp_add_in_reg_0_0; // @[FloatingPointDesigns.scala 1488:44]
  reg [23:0] cmpl_wire_temp_add_in_reg_0_1; // @[FloatingPointDesigns.scala 1488:44]
  wire [23:0] _cmpl_wire_temp_add_in_reg_0_0_T = ~wire_temp_add_in_reg_0_0; // @[FloatingPointDesigns.scala 1490:48]
  wire [23:0] _cmpl_wire_temp_add_in_reg_0_0_T_2 = 24'h1 + _cmpl_wire_temp_add_in_reg_0_0_T; // @[FloatingPointDesigns.scala 1490:46]
  wire [23:0] _cmpl_wire_temp_add_in_reg_0_1_T = ~wire_temp_add_in_reg_0_1; // @[FloatingPointDesigns.scala 1491:48]
  wire [23:0] _cmpl_wire_temp_add_in_reg_0_1_T_2 = 24'h1 + _cmpl_wire_temp_add_in_reg_0_1_T; // @[FloatingPointDesigns.scala 1491:46]
  wire [1:0] _adder_io_in_a_T = {sign_reg_4_1,sign_reg_4_0}; // @[FloatingPointDesigns.scala 1494:38]
  wire  _new_s_T = ~adder_io_out_c_reg_0; // @[FloatingPointDesigns.scala 1501:15]
  wire  new_s = ~adder_io_out_c_reg_0 & (sign_reg_5_0 | sign_reg_5_1) | sign_reg_5_0 & sign_reg_5_1; // @[FloatingPointDesigns.scala 1501:75]
  wire  _D_T_1 = sign_reg_5_0 ^ sign_reg_5_1; // @[FloatingPointDesigns.scala 1508:53]
  wire  D = _new_s_T | sign_reg_5_0 ^ sign_reg_5_1; // @[FloatingPointDesigns.scala 1508:35]
  wire  E = _new_s_T & ~adder_io_out_s_reg_0[23] | _new_s_T & ~_D_T_1 | adder_io_out_c_reg_0 & adder_io_out_s_reg_0[23]
     & _D_T_1; // @[FloatingPointDesigns.scala 1510:134]
  reg [23:0] cmpl_adder_io_out_s_reg_0; // @[FloatingPointDesigns.scala 1512:42]
  wire [23:0] _cmpl_adder_io_out_s_reg_0_T = ~adder_io_out_s_reg_1; // @[FloatingPointDesigns.scala 1515:43]
  wire [23:0] _cmpl_adder_io_out_s_reg_0_T_2 = 24'h1 + _cmpl_adder_io_out_s_reg_0_T; // @[FloatingPointDesigns.scala 1515:41]
  wire [1:0] _adder_result_T = {sign_reg_7_1,sign_reg_7_0}; // @[FloatingPointDesigns.scala 1519:53]
  wire [1:0] _leadingOne_T_25 = adder_result_reg_0[2] ? 2'h2 : {{1'd0}, adder_result_reg_0[1]}; // @[FloatingPointDesigns.scala 1522:70]
  wire [1:0] _leadingOne_T_26 = adder_result_reg_0[3] ? 2'h3 : _leadingOne_T_25; // @[FloatingPointDesigns.scala 1522:70]
  wire [2:0] _leadingOne_T_27 = adder_result_reg_0[4] ? 3'h4 : {{1'd0}, _leadingOne_T_26}; // @[FloatingPointDesigns.scala 1522:70]
  wire [2:0] _leadingOne_T_28 = adder_result_reg_0[5] ? 3'h5 : _leadingOne_T_27; // @[FloatingPointDesigns.scala 1522:70]
  wire [2:0] _leadingOne_T_29 = adder_result_reg_0[6] ? 3'h6 : _leadingOne_T_28; // @[FloatingPointDesigns.scala 1522:70]
  wire [2:0] _leadingOne_T_30 = adder_result_reg_0[7] ? 3'h7 : _leadingOne_T_29; // @[FloatingPointDesigns.scala 1522:70]
  wire [3:0] _leadingOne_T_31 = adder_result_reg_0[8] ? 4'h8 : {{1'd0}, _leadingOne_T_30}; // @[FloatingPointDesigns.scala 1522:70]
  wire [3:0] _leadingOne_T_32 = adder_result_reg_0[9] ? 4'h9 : _leadingOne_T_31; // @[FloatingPointDesigns.scala 1522:70]
  wire [3:0] _leadingOne_T_33 = adder_result_reg_0[10] ? 4'ha : _leadingOne_T_32; // @[FloatingPointDesigns.scala 1522:70]
  wire [3:0] _leadingOne_T_34 = adder_result_reg_0[11] ? 4'hb : _leadingOne_T_33; // @[FloatingPointDesigns.scala 1522:70]
  wire [3:0] _leadingOne_T_35 = adder_result_reg_0[12] ? 4'hc : _leadingOne_T_34; // @[FloatingPointDesigns.scala 1522:70]
  wire [3:0] _leadingOne_T_36 = adder_result_reg_0[13] ? 4'hd : _leadingOne_T_35; // @[FloatingPointDesigns.scala 1522:70]
  wire [3:0] _leadingOne_T_37 = adder_result_reg_0[14] ? 4'he : _leadingOne_T_36; // @[FloatingPointDesigns.scala 1522:70]
  wire [3:0] _leadingOne_T_38 = adder_result_reg_0[15] ? 4'hf : _leadingOne_T_37; // @[FloatingPointDesigns.scala 1522:70]
  wire [4:0] _leadingOne_T_39 = adder_result_reg_0[16] ? 5'h10 : {{1'd0}, _leadingOne_T_38}; // @[FloatingPointDesigns.scala 1522:70]
  wire [4:0] _leadingOne_T_40 = adder_result_reg_0[17] ? 5'h11 : _leadingOne_T_39; // @[FloatingPointDesigns.scala 1522:70]
  wire [4:0] _leadingOne_T_41 = adder_result_reg_0[18] ? 5'h12 : _leadingOne_T_40; // @[FloatingPointDesigns.scala 1522:70]
  wire [4:0] _leadingOne_T_42 = adder_result_reg_0[19] ? 5'h13 : _leadingOne_T_41; // @[FloatingPointDesigns.scala 1522:70]
  wire [4:0] _leadingOne_T_43 = adder_result_reg_0[20] ? 5'h14 : _leadingOne_T_42; // @[FloatingPointDesigns.scala 1522:70]
  wire [4:0] _leadingOne_T_44 = adder_result_reg_0[21] ? 5'h15 : _leadingOne_T_43; // @[FloatingPointDesigns.scala 1522:70]
  wire [4:0] _leadingOne_T_45 = adder_result_reg_0[22] ? 5'h16 : _leadingOne_T_44; // @[FloatingPointDesigns.scala 1522:70]
  wire [4:0] _leadingOne_T_46 = adder_result_reg_0[23] ? 5'h17 : _leadingOne_T_45; // @[FloatingPointDesigns.scala 1522:70]
  wire [5:0] leadingOne = _leadingOne_T_46 + 5'h1; // @[FloatingPointDesigns.scala 1522:77]
  wire [5:0] _subber2_io_in_b_T_1 = 6'h18 - leadingOne_reg_0; // @[FloatingPointDesigns.scala 1525:42]
  wire [7:0] exp_0 = _GEN_1[7:0]; // @[FloatingPointDesigns.scala 1387:19]
  wire [7:0] exp_1 = _GEN_3[7:0]; // @[FloatingPointDesigns.scala 1387:19]
  wire [7:0] _GEN_24 = subber_io_out_s; // @[FloatingPointDesigns.scala 1529:19 1538:27 1419:35]
  wire  _GEN_25 = subber_io_out_c; // @[FloatingPointDesigns.scala 1529:19 1539:27 1420:35]
  wire [23:0] _GEN_35 = adder_io_out_s; // @[FloatingPointDesigns.scala 1529:19 1554:29 1429:37]
  wire  _GEN_36 = adder_io_out_c; // @[FloatingPointDesigns.scala 1529:19 1555:29 1430:37]
  wire [7:0] _GEN_39 = subber2_io_out_s; // @[FloatingPointDesigns.scala 1529:19 1561:28 1445:36]
  wire  _GEN_40 = subber2_io_out_c; // @[FloatingPointDesigns.scala 1529:19 1562:28 1446:36]
  reg [31:0] reg_out_s; // @[FloatingPointDesigns.scala 1596:28]
  wire [8:0] _GEN_169 = {{1'd0}, ref_exp_reg_7}; // @[FloatingPointDesigns.scala 1613:29]
  wire [23:0] _new_out_frac_reg_0_T_2 = 24'h800000 - 24'h1; // @[FloatingPointDesigns.scala 1615:60]
  wire [7:0] _new_out_exp_reg_0_T_3 = ref_exp_reg_7 + 8'h1; // @[FloatingPointDesigns.scala 1617:48]
  wire [8:0] _GEN_142 = _GEN_169 == _T_2 ? _T_2 : {{1'd0}, _new_out_exp_reg_0_T_3}; // @[FloatingPointDesigns.scala 1613:66 1614:30 1617:30]
  wire [23:0] _GEN_143 = _GEN_169 == _T_2 ? _new_out_frac_reg_0_T_2 : {{1'd0}, adder_result_reg_2[23:1]}; // @[FloatingPointDesigns.scala 1613:66 1615:31 1618:31]
  wire [5:0] _new_out_frac_reg_0_T_6 = 6'h18 - leadingOne_reg_1; // @[FloatingPointDesigns.scala 1631:94]
  wire [85:0] _GEN_4 = {{63'd0}, adder_result_reg_2[22:0]}; // @[FloatingPointDesigns.scala 1631:73]
  wire [85:0] _new_out_frac_reg_0_T_7 = _GEN_4 << _new_out_frac_reg_0_T_6; // @[FloatingPointDesigns.scala 1631:73]
  wire [7:0] _GEN_144 = subber2_out_c_reg_0 ? 8'h1 : subber2_out_s_reg_0; // @[FloatingPointDesigns.scala 1626:46 1627:32 1630:32]
  wire [85:0] _GEN_145 = subber2_out_c_reg_0 ? 86'h0 : _new_out_frac_reg_0_T_7; // @[FloatingPointDesigns.scala 1626:46 1628:33 1631:33]
  wire [7:0] _GEN_146 = leadingOne_reg_1 == 6'h1 & adder_result_reg_2 == 24'h0 & ((sign_reg_10_0 ^ sign_reg_10_1) &
    io_in_a_reg_10[30:0] == io_in_b_reg_10[30:0]) ? 8'h0 : _GEN_144; // @[FloatingPointDesigns.scala 1622:184 1623:30]
  wire [85:0] _GEN_147 = leadingOne_reg_1 == 6'h1 & adder_result_reg_2 == 24'h0 & ((sign_reg_10_0 ^ sign_reg_10_1) &
    io_in_a_reg_10[30:0] == io_in_b_reg_10[30:0]) ? 86'h0 : _GEN_145; // @[FloatingPointDesigns.scala 1622:184 1624:31]
  wire  _GEN_148 = D_reg_4 ? new_s_reg_4 : new_s_reg_5; // @[FloatingPointDesigns.scala 1620:36 1621:22 1432:35]
  wire [7:0] _GEN_149 = D_reg_4 ? _GEN_146 : new_out_exp_reg_0; // @[FloatingPointDesigns.scala 1434:35 1620:36]
  wire [85:0] _GEN_150 = D_reg_4 ? _GEN_147 : {{63'd0}, new_out_frac_reg_0}; // @[FloatingPointDesigns.scala 1433:35 1620:36]
  wire  _GEN_151 = ~D_reg_4 ? new_s_reg_4 : _GEN_148; // @[FloatingPointDesigns.scala 1611:36 1612:22]
  wire [8:0] _GEN_152 = ~D_reg_4 ? _GEN_142 : {{1'd0}, _GEN_149}; // @[FloatingPointDesigns.scala 1611:36]
  wire [85:0] _GEN_153 = ~D_reg_4 ? {{62'd0}, _GEN_143} : _GEN_150; // @[FloatingPointDesigns.scala 1611:36]
  wire [8:0] _GEN_155 = E_reg_4 ? {{1'd0}, ref_exp_reg_7} : _GEN_152; // @[FloatingPointDesigns.scala 1607:36 1609:28]
  wire [85:0] _GEN_156 = E_reg_4 ? {{63'd0}, adder_result_reg_2[22:0]} : _GEN_153; // @[FloatingPointDesigns.scala 1607:36 1610:29]
  wire [85:0] _GEN_158 = sub_exp_reg_7 >= 8'h17 ? {{63'd0}, ref_frac_reg_7} : _GEN_156; // @[FloatingPointDesigns.scala 1603:48 1605:29]
  wire [8:0] _GEN_159 = sub_exp_reg_7 >= 8'h17 ? {{1'd0}, ref_exp_reg_7} : _GEN_155; // @[FloatingPointDesigns.scala 1603:48 1606:28]
  wire [8:0] _GEN_161 = io_in_a_reg_10[30:0] == 31'h0 & io_in_b_reg_10[30:0] == 31'h0 ? 9'h0 : _GEN_159; // @[FloatingPointDesigns.scala 1599:86 1601:28]
  wire [85:0] _GEN_162 = io_in_a_reg_10[30:0] == 31'h0 & io_in_b_reg_10[30:0] == 31'h0 ? 86'h0 : _GEN_158; // @[FloatingPointDesigns.scala 1599:86 1602:29]
  wire [31:0] _reg_out_s_T_1 = {new_s_reg_5,new_out_exp_reg_0,new_out_frac_reg_0}; // @[FloatingPointDesigns.scala 1635:55]
  wire [85:0] _GEN_170 = reset ? 86'h0 : _GEN_162; // @[FloatingPointDesigns.scala 1433:{35,35}]
  wire [8:0] _GEN_171 = reset ? 9'h0 : _GEN_161; // @[FloatingPointDesigns.scala 1434:{35,35}]
  full_subber subber ( // @[FloatingPointDesigns.scala 1456:24]
    .io_in_a(subber_io_in_a),
    .io_in_b(subber_io_in_b),
    .io_out_s(subber_io_out_s),
    .io_out_c(subber_io_out_c)
  );
  full_adder_128 adder ( // @[FloatingPointDesigns.scala 1462:23]
    .io_in_a(adder_io_in_a),
    .io_in_b(adder_io_in_b),
    .io_out_s(adder_io_out_s),
    .io_out_c(adder_io_out_c)
  );
  full_subber subber2 ( // @[FloatingPointDesigns.scala 1523:25]
    .io_in_a(subber2_io_in_a),
    .io_in_b(subber2_io_in_b),
    .io_out_s(subber2_io_out_s),
    .io_out_c(subber2_io_out_c)
  );
  assign io_out_s = reg_out_s; // @[FloatingPointDesigns.scala 1597:14]
  assign subber_io_in_a = exp_reg_0_0; // @[FloatingPointDesigns.scala 1457:20]
  assign subber_io_in_b = exp_reg_0_1; // @[FloatingPointDesigns.scala 1458:20]
  assign adder_io_in_a = _adder_io_in_a_T == 2'h1 ? cmpl_wire_temp_add_in_reg_0_0 : wire_temp_add_in_reg_1_0; // @[FloatingPointDesigns.scala 1494:25]
  assign adder_io_in_b = _adder_io_in_a_T == 2'h2 ? cmpl_wire_temp_add_in_reg_0_1 : wire_temp_add_in_reg_1_1; // @[FloatingPointDesigns.scala 1495:25]
  assign subber2_io_in_a = ref_exp_reg_6; // @[FloatingPointDesigns.scala 1524:21]
  assign subber2_io_in_b = {{2'd0}, _subber2_io_in_b_T_1}; // @[FloatingPointDesigns.scala 1525:21]
  always @(posedge clock) begin
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_0_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_0_0 <= sign_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_0_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_0_1 <= sign_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_1_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_1_0 <= sign_reg_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_1_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_1_1 <= sign_reg_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_2_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_2_0 <= sign_reg_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_2_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_2_1 <= sign_reg_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_3_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_3_0 <= sign_reg_2_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_3_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_3_1 <= sign_reg_2_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_4_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_4_0 <= sign_reg_3_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_4_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_4_1 <= sign_reg_3_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_5_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_5_0 <= sign_reg_4_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_5_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_5_1 <= sign_reg_4_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_6_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_6_0 <= sign_reg_5_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_6_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_6_1 <= sign_reg_5_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_7_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_7_0 <= sign_reg_6_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_7_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_7_1 <= sign_reg_6_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_8_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_8_0 <= sign_reg_7_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_8_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_8_1 <= sign_reg_7_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_9_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_9_0 <= sign_reg_8_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_9_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_9_1 <= sign_reg_8_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_10_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_10_0 <= sign_reg_9_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_10_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_10_1 <= sign_reg_9_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1415:28]
      exp_reg_0_0 <= 8'h0; // @[FloatingPointDesigns.scala 1415:28]
    end else begin
      exp_reg_0_0 <= exp_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1415:28]
      exp_reg_0_1 <= 8'h0; // @[FloatingPointDesigns.scala 1415:28]
    end else begin
      exp_reg_0_1 <= exp_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1415:28]
      exp_reg_1_0 <= 8'h0; // @[FloatingPointDesigns.scala 1415:28]
    end else begin
      exp_reg_1_0 <= exp_reg_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1415:28]
      exp_reg_1_1 <= 8'h0; // @[FloatingPointDesigns.scala 1415:28]
    end else begin
      exp_reg_1_1 <= exp_reg_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1415:28]
      exp_reg_2_0 <= 8'h0; // @[FloatingPointDesigns.scala 1415:28]
    end else begin
      exp_reg_2_0 <= exp_reg_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1415:28]
      exp_reg_2_1 <= 8'h0; // @[FloatingPointDesigns.scala 1415:28]
    end else begin
      exp_reg_2_1 <= exp_reg_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1416:28]
      frac_reg_0_0 <= 23'h0; // @[FloatingPointDesigns.scala 1416:28]
    end else begin
      frac_reg_0_0 <= frac_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1416:28]
      frac_reg_0_1 <= 23'h0; // @[FloatingPointDesigns.scala 1416:28]
    end else begin
      frac_reg_0_1 <= frac_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1416:28]
      frac_reg_1_0 <= 23'h0; // @[FloatingPointDesigns.scala 1416:28]
    end else begin
      frac_reg_1_0 <= frac_reg_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1416:28]
      frac_reg_1_1 <= 23'h0; // @[FloatingPointDesigns.scala 1416:28]
    end else begin
      frac_reg_1_1 <= frac_reg_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1416:28]
      frac_reg_2_0 <= 23'h0; // @[FloatingPointDesigns.scala 1416:28]
    end else begin
      frac_reg_2_0 <= frac_reg_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1416:28]
      frac_reg_2_1 <= 23'h0; // @[FloatingPointDesigns.scala 1416:28]
    end else begin
      frac_reg_2_1 <= frac_reg_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1417:28]
      wfrac_reg_0_0 <= 24'h0; // @[FloatingPointDesigns.scala 1417:28]
    end else begin
      wfrac_reg_0_0 <= whole_frac_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1417:28]
      wfrac_reg_0_1 <= 24'h0; // @[FloatingPointDesigns.scala 1417:28]
    end else begin
      wfrac_reg_0_1 <= whole_frac_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1417:28]
      wfrac_reg_1_0 <= 24'h0; // @[FloatingPointDesigns.scala 1417:28]
    end else begin
      wfrac_reg_1_0 <= wfrac_reg_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1417:28]
      wfrac_reg_1_1 <= 24'h0; // @[FloatingPointDesigns.scala 1417:28]
    end else begin
      wfrac_reg_1_1 <= wfrac_reg_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1417:28]
      wfrac_reg_2_0 <= 24'h0; // @[FloatingPointDesigns.scala 1417:28]
    end else begin
      wfrac_reg_2_0 <= wfrac_reg_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1417:28]
      wfrac_reg_2_1 <= 24'h0; // @[FloatingPointDesigns.scala 1417:28]
    end else begin
      wfrac_reg_2_1 <= wfrac_reg_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1419:35]
      subber_out_s_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1419:35]
    end else begin
      subber_out_s_reg_0 <= _GEN_24;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1419:35]
      subber_out_s_reg_1 <= 8'h0; // @[FloatingPointDesigns.scala 1419:35]
    end else begin
      subber_out_s_reg_1 <= subber_out_s_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1420:35]
      subber_out_c_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1420:35]
    end else begin
      subber_out_c_reg_0 <= _GEN_25;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1420:35]
      subber_out_c_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1420:35]
    end else begin
      subber_out_c_reg_1 <= subber_out_c_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1422:39]
      wire_temp_add_in_reg_0_0 <= 24'h0; // @[FloatingPointDesigns.scala 1422:39]
    end else if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1472:39]
      wire_temp_add_in_reg_0_0 <= _wire_temp_add_in_0_T; // @[FloatingPointDesigns.scala 1477:27]
    end else begin
      wire_temp_add_in_reg_0_0 <= wfrac_reg_2_0; // @[FloatingPointDesigns.scala 1484:27]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1422:39]
      wire_temp_add_in_reg_0_1 <= 24'h0; // @[FloatingPointDesigns.scala 1422:39]
    end else if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1472:39]
      wire_temp_add_in_reg_0_1 <= wfrac_reg_2_1; // @[FloatingPointDesigns.scala 1478:27]
    end else begin
      wire_temp_add_in_reg_0_1 <= _wire_temp_add_in_1_T; // @[FloatingPointDesigns.scala 1485:27]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1422:39]
      wire_temp_add_in_reg_1_0 <= 24'h0; // @[FloatingPointDesigns.scala 1422:39]
    end else begin
      wire_temp_add_in_reg_1_0 <= wire_temp_add_in_reg_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1422:39]
      wire_temp_add_in_reg_1_1 <= 24'h0; // @[FloatingPointDesigns.scala 1422:39]
    end else begin
      wire_temp_add_in_reg_1_1 <= wire_temp_add_in_reg_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1424:31]
      ref_s_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1424:31]
    end else if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1472:39]
      ref_s_reg_0 <= sign_reg_2_1; // @[FloatingPointDesigns.scala 1475:13]
    end else begin
      ref_s_reg_0 <= sign_reg_2_0; // @[FloatingPointDesigns.scala 1482:13]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1424:31]
      ref_s_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1424:31]
    end else begin
      ref_s_reg_1 <= ref_s_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1424:31]
      ref_s_reg_2 <= 1'h0; // @[FloatingPointDesigns.scala 1424:31]
    end else begin
      ref_s_reg_2 <= ref_s_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1424:31]
      ref_s_reg_3 <= 1'h0; // @[FloatingPointDesigns.scala 1424:31]
    end else begin
      ref_s_reg_3 <= ref_s_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1424:31]
      ref_s_reg_4 <= 1'h0; // @[FloatingPointDesigns.scala 1424:31]
    end else begin
      ref_s_reg_4 <= ref_s_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1424:31]
      ref_s_reg_5 <= 1'h0; // @[FloatingPointDesigns.scala 1424:31]
    end else begin
      ref_s_reg_5 <= ref_s_reg_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1424:31]
      ref_s_reg_6 <= 1'h0; // @[FloatingPointDesigns.scala 1424:31]
    end else begin
      ref_s_reg_6 <= ref_s_reg_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1424:31]
      ref_s_reg_7 <= 1'h0; // @[FloatingPointDesigns.scala 1424:31]
    end else begin
      ref_s_reg_7 <= ref_s_reg_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1425:31]
      ref_frac_reg_0 <= 23'h0; // @[FloatingPointDesigns.scala 1425:31]
    end else if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1472:39]
      ref_frac_reg_0 <= frac_reg_2_1; // @[FloatingPointDesigns.scala 1476:16]
    end else begin
      ref_frac_reg_0 <= frac_reg_2_0; // @[FloatingPointDesigns.scala 1483:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1425:31]
      ref_frac_reg_1 <= 23'h0; // @[FloatingPointDesigns.scala 1425:31]
    end else begin
      ref_frac_reg_1 <= ref_frac_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1425:31]
      ref_frac_reg_2 <= 23'h0; // @[FloatingPointDesigns.scala 1425:31]
    end else begin
      ref_frac_reg_2 <= ref_frac_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1425:31]
      ref_frac_reg_3 <= 23'h0; // @[FloatingPointDesigns.scala 1425:31]
    end else begin
      ref_frac_reg_3 <= ref_frac_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1425:31]
      ref_frac_reg_4 <= 23'h0; // @[FloatingPointDesigns.scala 1425:31]
    end else begin
      ref_frac_reg_4 <= ref_frac_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1425:31]
      ref_frac_reg_5 <= 23'h0; // @[FloatingPointDesigns.scala 1425:31]
    end else begin
      ref_frac_reg_5 <= ref_frac_reg_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1425:31]
      ref_frac_reg_6 <= 23'h0; // @[FloatingPointDesigns.scala 1425:31]
    end else begin
      ref_frac_reg_6 <= ref_frac_reg_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1425:31]
      ref_frac_reg_7 <= 23'h0; // @[FloatingPointDesigns.scala 1425:31]
    end else begin
      ref_frac_reg_7 <= ref_frac_reg_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1426:31]
      ref_exp_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1426:31]
    end else if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1472:39]
      ref_exp_reg_0 <= exp_reg_2_1; // @[FloatingPointDesigns.scala 1473:15]
    end else begin
      ref_exp_reg_0 <= exp_reg_2_0; // @[FloatingPointDesigns.scala 1480:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1426:31]
      ref_exp_reg_1 <= 8'h0; // @[FloatingPointDesigns.scala 1426:31]
    end else begin
      ref_exp_reg_1 <= ref_exp_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1426:31]
      ref_exp_reg_2 <= 8'h0; // @[FloatingPointDesigns.scala 1426:31]
    end else begin
      ref_exp_reg_2 <= ref_exp_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1426:31]
      ref_exp_reg_3 <= 8'h0; // @[FloatingPointDesigns.scala 1426:31]
    end else begin
      ref_exp_reg_3 <= ref_exp_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1426:31]
      ref_exp_reg_4 <= 8'h0; // @[FloatingPointDesigns.scala 1426:31]
    end else begin
      ref_exp_reg_4 <= ref_exp_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1426:31]
      ref_exp_reg_5 <= 8'h0; // @[FloatingPointDesigns.scala 1426:31]
    end else begin
      ref_exp_reg_5 <= ref_exp_reg_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1426:31]
      ref_exp_reg_6 <= 8'h0; // @[FloatingPointDesigns.scala 1426:31]
    end else begin
      ref_exp_reg_6 <= ref_exp_reg_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1426:31]
      ref_exp_reg_7 <= 8'h0; // @[FloatingPointDesigns.scala 1426:31]
    end else begin
      ref_exp_reg_7 <= ref_exp_reg_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1427:31]
      sub_exp_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1427:31]
    end else if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1472:39]
      sub_exp_reg_0 <= cmpl_subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1474:15]
    end else begin
      sub_exp_reg_0 <= subber_out_s_reg_1; // @[FloatingPointDesigns.scala 1481:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1427:31]
      sub_exp_reg_1 <= 8'h0; // @[FloatingPointDesigns.scala 1427:31]
    end else begin
      sub_exp_reg_1 <= sub_exp_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1427:31]
      sub_exp_reg_2 <= 8'h0; // @[FloatingPointDesigns.scala 1427:31]
    end else begin
      sub_exp_reg_2 <= sub_exp_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1427:31]
      sub_exp_reg_3 <= 8'h0; // @[FloatingPointDesigns.scala 1427:31]
    end else begin
      sub_exp_reg_3 <= sub_exp_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1427:31]
      sub_exp_reg_4 <= 8'h0; // @[FloatingPointDesigns.scala 1427:31]
    end else begin
      sub_exp_reg_4 <= sub_exp_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1427:31]
      sub_exp_reg_5 <= 8'h0; // @[FloatingPointDesigns.scala 1427:31]
    end else begin
      sub_exp_reg_5 <= sub_exp_reg_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1427:31]
      sub_exp_reg_6 <= 8'h0; // @[FloatingPointDesigns.scala 1427:31]
    end else begin
      sub_exp_reg_6 <= sub_exp_reg_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1427:31]
      sub_exp_reg_7 <= 8'h0; // @[FloatingPointDesigns.scala 1427:31]
    end else begin
      sub_exp_reg_7 <= sub_exp_reg_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1429:37]
      adder_io_out_s_reg_0 <= 24'h0; // @[FloatingPointDesigns.scala 1429:37]
    end else begin
      adder_io_out_s_reg_0 <= _GEN_35;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1429:37]
      adder_io_out_s_reg_1 <= 24'h0; // @[FloatingPointDesigns.scala 1429:37]
    end else begin
      adder_io_out_s_reg_1 <= adder_io_out_s_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1429:37]
      adder_io_out_s_reg_2 <= 24'h0; // @[FloatingPointDesigns.scala 1429:37]
    end else begin
      adder_io_out_s_reg_2 <= adder_io_out_s_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1430:37]
      adder_io_out_c_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1430:37]
    end else begin
      adder_io_out_c_reg_0 <= _GEN_36;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1432:35]
      new_s_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1432:35]
    end else begin
      new_s_reg_0 <= new_s;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1432:35]
      new_s_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1432:35]
    end else begin
      new_s_reg_1 <= new_s_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1432:35]
      new_s_reg_2 <= 1'h0; // @[FloatingPointDesigns.scala 1432:35]
    end else begin
      new_s_reg_2 <= new_s_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1432:35]
      new_s_reg_3 <= 1'h0; // @[FloatingPointDesigns.scala 1432:35]
    end else begin
      new_s_reg_3 <= new_s_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1432:35]
      new_s_reg_4 <= 1'h0; // @[FloatingPointDesigns.scala 1432:35]
    end else begin
      new_s_reg_4 <= new_s_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1432:35]
      new_s_reg_5 <= 1'h0; // @[FloatingPointDesigns.scala 1432:35]
    end else if (io_in_a_reg_10[30:0] == 31'h0 & io_in_b_reg_10[30:0] == 31'h0) begin // @[FloatingPointDesigns.scala 1599:86]
      new_s_reg_5 <= 1'h0; // @[FloatingPointDesigns.scala 1600:22]
    end else if (sub_exp_reg_7 >= 8'h17) begin // @[FloatingPointDesigns.scala 1603:48]
      new_s_reg_5 <= ref_s_reg_7; // @[FloatingPointDesigns.scala 1604:22]
    end else if (E_reg_4) begin // @[FloatingPointDesigns.scala 1607:36]
      new_s_reg_5 <= new_s_reg_4; // @[FloatingPointDesigns.scala 1608:22]
    end else begin
      new_s_reg_5 <= _GEN_151;
    end
    new_out_frac_reg_0 <= _GEN_170[22:0]; // @[FloatingPointDesigns.scala 1433:{35,35}]
    new_out_exp_reg_0 <= _GEN_171[7:0]; // @[FloatingPointDesigns.scala 1434:{35,35}]
    if (reset) begin // @[FloatingPointDesigns.scala 1435:24]
      E_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1435:24]
    end else begin
      E_reg_0 <= E;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1435:24]
      E_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1435:24]
    end else begin
      E_reg_1 <= E_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1435:24]
      E_reg_2 <= 1'h0; // @[FloatingPointDesigns.scala 1435:24]
    end else begin
      E_reg_2 <= E_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1435:24]
      E_reg_3 <= 1'h0; // @[FloatingPointDesigns.scala 1435:24]
    end else begin
      E_reg_3 <= E_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1435:24]
      E_reg_4 <= 1'h0; // @[FloatingPointDesigns.scala 1435:24]
    end else begin
      E_reg_4 <= E_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1436:24]
      D_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1436:24]
    end else begin
      D_reg_0 <= D;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1436:24]
      D_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1436:24]
    end else begin
      D_reg_1 <= D_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1436:24]
      D_reg_2 <= 1'h0; // @[FloatingPointDesigns.scala 1436:24]
    end else begin
      D_reg_2 <= D_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1436:24]
      D_reg_3 <= 1'h0; // @[FloatingPointDesigns.scala 1436:24]
    end else begin
      D_reg_3 <= D_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1436:24]
      D_reg_4 <= 1'h0; // @[FloatingPointDesigns.scala 1436:24]
    end else begin
      D_reg_4 <= D_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1438:35]
      adder_result_reg_0 <= 24'h0; // @[FloatingPointDesigns.scala 1438:35]
    end else if (new_s_reg_1 & ^_adder_result_T) begin // @[FloatingPointDesigns.scala 1519:24]
      adder_result_reg_0 <= cmpl_adder_io_out_s_reg_0;
    end else begin
      adder_result_reg_0 <= adder_io_out_s_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1438:35]
      adder_result_reg_1 <= 24'h0; // @[FloatingPointDesigns.scala 1438:35]
    end else begin
      adder_result_reg_1 <= adder_result_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1438:35]
      adder_result_reg_2 <= 24'h0; // @[FloatingPointDesigns.scala 1438:35]
    end else begin
      adder_result_reg_2 <= adder_result_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1440:33]
      leadingOne_reg_0 <= 6'h0; // @[FloatingPointDesigns.scala 1440:33]
    end else begin
      leadingOne_reg_0 <= leadingOne;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1440:33]
      leadingOne_reg_1 <= 6'h0; // @[FloatingPointDesigns.scala 1440:33]
    end else begin
      leadingOne_reg_1 <= leadingOne_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_0 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_0 <= io_in_a;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_1 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_1 <= io_in_a_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_2 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_2 <= io_in_a_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_3 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_3 <= io_in_a_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_4 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_4 <= io_in_a_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_5 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_5 <= io_in_a_reg_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_6 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_6 <= io_in_a_reg_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_7 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_7 <= io_in_a_reg_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_8 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_8 <= io_in_a_reg_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_9 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_9 <= io_in_a_reg_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_10 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_10 <= io_in_a_reg_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_0 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_0 <= io_in_b;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_1 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_1 <= io_in_b_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_2 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_2 <= io_in_b_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_3 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_3 <= io_in_b_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_4 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_4 <= io_in_b_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_5 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_5 <= io_in_b_reg_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_6 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_6 <= io_in_b_reg_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_7 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_7 <= io_in_b_reg_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_8 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_8 <= io_in_b_reg_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_9 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_9 <= io_in_b_reg_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_10 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_10 <= io_in_b_reg_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1445:36]
      subber2_out_s_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1445:36]
    end else begin
      subber2_out_s_reg_0 <= _GEN_39;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1446:36]
      subber2_out_c_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1446:36]
    end else begin
      subber2_out_c_reg_0 <= _GEN_40;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1467:40]
      cmpl_subber_out_s_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1467:40]
    end else begin
      cmpl_subber_out_s_reg_0 <= _cmpl_subber_out_s_reg_0_T_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1488:44]
      cmpl_wire_temp_add_in_reg_0_0 <= 24'h0; // @[FloatingPointDesigns.scala 1488:44]
    end else begin
      cmpl_wire_temp_add_in_reg_0_0 <= _cmpl_wire_temp_add_in_reg_0_0_T_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1488:44]
      cmpl_wire_temp_add_in_reg_0_1 <= 24'h0; // @[FloatingPointDesigns.scala 1488:44]
    end else begin
      cmpl_wire_temp_add_in_reg_0_1 <= _cmpl_wire_temp_add_in_reg_0_1_T_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1512:42]
      cmpl_adder_io_out_s_reg_0 <= 24'h0; // @[FloatingPointDesigns.scala 1512:42]
    end else begin
      cmpl_adder_io_out_s_reg_0 <= _cmpl_adder_io_out_s_reg_0_T_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1596:28]
      reg_out_s <= 32'h0; // @[FloatingPointDesigns.scala 1596:28]
    end else begin
      reg_out_s <= _reg_out_s_T_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sign_reg_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sign_reg_0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sign_reg_1_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  sign_reg_1_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  sign_reg_2_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  sign_reg_2_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  sign_reg_3_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  sign_reg_3_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  sign_reg_4_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sign_reg_4_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  sign_reg_5_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  sign_reg_5_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  sign_reg_6_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  sign_reg_6_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  sign_reg_7_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  sign_reg_7_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  sign_reg_8_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  sign_reg_8_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  sign_reg_9_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sign_reg_9_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  sign_reg_10_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  sign_reg_10_1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  exp_reg_0_0 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  exp_reg_0_1 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  exp_reg_1_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  exp_reg_1_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  exp_reg_2_0 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  exp_reg_2_1 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  frac_reg_0_0 = _RAND_28[22:0];
  _RAND_29 = {1{`RANDOM}};
  frac_reg_0_1 = _RAND_29[22:0];
  _RAND_30 = {1{`RANDOM}};
  frac_reg_1_0 = _RAND_30[22:0];
  _RAND_31 = {1{`RANDOM}};
  frac_reg_1_1 = _RAND_31[22:0];
  _RAND_32 = {1{`RANDOM}};
  frac_reg_2_0 = _RAND_32[22:0];
  _RAND_33 = {1{`RANDOM}};
  frac_reg_2_1 = _RAND_33[22:0];
  _RAND_34 = {1{`RANDOM}};
  wfrac_reg_0_0 = _RAND_34[23:0];
  _RAND_35 = {1{`RANDOM}};
  wfrac_reg_0_1 = _RAND_35[23:0];
  _RAND_36 = {1{`RANDOM}};
  wfrac_reg_1_0 = _RAND_36[23:0];
  _RAND_37 = {1{`RANDOM}};
  wfrac_reg_1_1 = _RAND_37[23:0];
  _RAND_38 = {1{`RANDOM}};
  wfrac_reg_2_0 = _RAND_38[23:0];
  _RAND_39 = {1{`RANDOM}};
  wfrac_reg_2_1 = _RAND_39[23:0];
  _RAND_40 = {1{`RANDOM}};
  subber_out_s_reg_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  subber_out_s_reg_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  subber_out_c_reg_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  subber_out_c_reg_1 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  wire_temp_add_in_reg_0_0 = _RAND_44[23:0];
  _RAND_45 = {1{`RANDOM}};
  wire_temp_add_in_reg_0_1 = _RAND_45[23:0];
  _RAND_46 = {1{`RANDOM}};
  wire_temp_add_in_reg_1_0 = _RAND_46[23:0];
  _RAND_47 = {1{`RANDOM}};
  wire_temp_add_in_reg_1_1 = _RAND_47[23:0];
  _RAND_48 = {1{`RANDOM}};
  ref_s_reg_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  ref_s_reg_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  ref_s_reg_2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  ref_s_reg_3 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  ref_s_reg_4 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  ref_s_reg_5 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  ref_s_reg_6 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  ref_s_reg_7 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  ref_frac_reg_0 = _RAND_56[22:0];
  _RAND_57 = {1{`RANDOM}};
  ref_frac_reg_1 = _RAND_57[22:0];
  _RAND_58 = {1{`RANDOM}};
  ref_frac_reg_2 = _RAND_58[22:0];
  _RAND_59 = {1{`RANDOM}};
  ref_frac_reg_3 = _RAND_59[22:0];
  _RAND_60 = {1{`RANDOM}};
  ref_frac_reg_4 = _RAND_60[22:0];
  _RAND_61 = {1{`RANDOM}};
  ref_frac_reg_5 = _RAND_61[22:0];
  _RAND_62 = {1{`RANDOM}};
  ref_frac_reg_6 = _RAND_62[22:0];
  _RAND_63 = {1{`RANDOM}};
  ref_frac_reg_7 = _RAND_63[22:0];
  _RAND_64 = {1{`RANDOM}};
  ref_exp_reg_0 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  ref_exp_reg_1 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  ref_exp_reg_2 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  ref_exp_reg_3 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  ref_exp_reg_4 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  ref_exp_reg_5 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  ref_exp_reg_6 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  ref_exp_reg_7 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  sub_exp_reg_0 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  sub_exp_reg_1 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  sub_exp_reg_2 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  sub_exp_reg_3 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  sub_exp_reg_4 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  sub_exp_reg_5 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  sub_exp_reg_6 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  sub_exp_reg_7 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  adder_io_out_s_reg_0 = _RAND_80[23:0];
  _RAND_81 = {1{`RANDOM}};
  adder_io_out_s_reg_1 = _RAND_81[23:0];
  _RAND_82 = {1{`RANDOM}};
  adder_io_out_s_reg_2 = _RAND_82[23:0];
  _RAND_83 = {1{`RANDOM}};
  adder_io_out_c_reg_0 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  new_s_reg_0 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  new_s_reg_1 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  new_s_reg_2 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  new_s_reg_3 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  new_s_reg_4 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  new_s_reg_5 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  new_out_frac_reg_0 = _RAND_90[22:0];
  _RAND_91 = {1{`RANDOM}};
  new_out_exp_reg_0 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  E_reg_0 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  E_reg_1 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  E_reg_2 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  E_reg_3 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  E_reg_4 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  D_reg_0 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  D_reg_1 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  D_reg_2 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  D_reg_3 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  D_reg_4 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  adder_result_reg_0 = _RAND_102[23:0];
  _RAND_103 = {1{`RANDOM}};
  adder_result_reg_1 = _RAND_103[23:0];
  _RAND_104 = {1{`RANDOM}};
  adder_result_reg_2 = _RAND_104[23:0];
  _RAND_105 = {1{`RANDOM}};
  leadingOne_reg_0 = _RAND_105[5:0];
  _RAND_106 = {1{`RANDOM}};
  leadingOne_reg_1 = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  io_in_a_reg_0 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  io_in_a_reg_1 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  io_in_a_reg_2 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  io_in_a_reg_3 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  io_in_a_reg_4 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  io_in_a_reg_5 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  io_in_a_reg_6 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  io_in_a_reg_7 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  io_in_a_reg_8 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  io_in_a_reg_9 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  io_in_a_reg_10 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  io_in_b_reg_0 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  io_in_b_reg_1 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  io_in_b_reg_2 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  io_in_b_reg_3 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  io_in_b_reg_4 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  io_in_b_reg_5 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  io_in_b_reg_6 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  io_in_b_reg_7 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  io_in_b_reg_8 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  io_in_b_reg_9 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  io_in_b_reg_10 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  subber2_out_s_reg_0 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  subber2_out_c_reg_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  cmpl_subber_out_s_reg_0 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  cmpl_wire_temp_add_in_reg_0_0 = _RAND_132[23:0];
  _RAND_133 = {1{`RANDOM}};
  cmpl_wire_temp_add_in_reg_0_1 = _RAND_133[23:0];
  _RAND_134 = {1{`RANDOM}};
  cmpl_adder_io_out_s_reg_0 = _RAND_134[23:0];
  _RAND_135 = {1{`RANDOM}};
  reg_out_s = _RAND_135[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FP_DDOT_dp(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_0,
  input  [31:0] io_in_a_1,
  input  [31:0] io_in_a_2,
  input  [31:0] io_in_a_3,
  input  [31:0] io_in_a_4,
  input  [31:0] io_in_a_5,
  input  [31:0] io_in_a_6,
  input  [31:0] io_in_a_7,
  input  [31:0] io_in_a_8,
  input  [31:0] io_in_a_9,
  input  [31:0] io_in_a_10,
  input  [31:0] io_in_a_11,
  input  [31:0] io_in_a_12,
  input  [31:0] io_in_a_13,
  input  [31:0] io_in_a_14,
  input  [31:0] io_in_a_15,
  input  [31:0] io_in_a_16,
  input  [31:0] io_in_a_17,
  input  [31:0] io_in_a_18,
  input  [31:0] io_in_a_19,
  input  [31:0] io_in_a_20,
  input  [31:0] io_in_a_21,
  input  [31:0] io_in_a_22,
  input  [31:0] io_in_a_23,
  input  [31:0] io_in_a_24,
  input  [31:0] io_in_a_25,
  input  [31:0] io_in_a_26,
  input  [31:0] io_in_a_27,
  input  [31:0] io_in_a_28,
  input  [31:0] io_in_a_29,
  input  [31:0] io_in_a_30,
  input  [31:0] io_in_a_31,
  input  [31:0] io_in_a_32,
  input  [31:0] io_in_a_33,
  input  [31:0] io_in_a_34,
  input  [31:0] io_in_a_35,
  input  [31:0] io_in_a_36,
  input  [31:0] io_in_a_37,
  input  [31:0] io_in_a_38,
  input  [31:0] io_in_a_39,
  input  [31:0] io_in_a_40,
  input  [31:0] io_in_a_41,
  input  [31:0] io_in_a_42,
  input  [31:0] io_in_a_43,
  input  [31:0] io_in_a_44,
  input  [31:0] io_in_a_45,
  input  [31:0] io_in_a_46,
  input  [31:0] io_in_a_47,
  input  [31:0] io_in_a_48,
  input  [31:0] io_in_a_49,
  input  [31:0] io_in_a_50,
  input  [31:0] io_in_a_51,
  input  [31:0] io_in_a_52,
  input  [31:0] io_in_a_53,
  input  [31:0] io_in_a_54,
  input  [31:0] io_in_a_55,
  input  [31:0] io_in_a_56,
  input  [31:0] io_in_a_57,
  input  [31:0] io_in_a_58,
  input  [31:0] io_in_a_59,
  input  [31:0] io_in_a_60,
  input  [31:0] io_in_a_61,
  input  [31:0] io_in_a_62,
  input  [31:0] io_in_a_63,
  input  [31:0] io_in_a_64,
  input  [31:0] io_in_a_65,
  input  [31:0] io_in_a_66,
  input  [31:0] io_in_a_67,
  input  [31:0] io_in_a_68,
  input  [31:0] io_in_a_69,
  input  [31:0] io_in_a_70,
  input  [31:0] io_in_a_71,
  input  [31:0] io_in_a_72,
  input  [31:0] io_in_a_73,
  input  [31:0] io_in_a_74,
  input  [31:0] io_in_a_75,
  input  [31:0] io_in_a_76,
  input  [31:0] io_in_a_77,
  input  [31:0] io_in_a_78,
  input  [31:0] io_in_a_79,
  input  [31:0] io_in_a_80,
  input  [31:0] io_in_a_81,
  input  [31:0] io_in_a_82,
  input  [31:0] io_in_a_83,
  input  [31:0] io_in_a_84,
  input  [31:0] io_in_a_85,
  input  [31:0] io_in_a_86,
  input  [31:0] io_in_a_87,
  input  [31:0] io_in_a_88,
  input  [31:0] io_in_a_89,
  input  [31:0] io_in_a_90,
  input  [31:0] io_in_a_91,
  input  [31:0] io_in_a_92,
  input  [31:0] io_in_a_93,
  input  [31:0] io_in_a_94,
  input  [31:0] io_in_a_95,
  input  [31:0] io_in_a_96,
  input  [31:0] io_in_a_97,
  input  [31:0] io_in_a_98,
  input  [31:0] io_in_a_99,
  input  [31:0] io_in_a_100,
  input  [31:0] io_in_a_101,
  input  [31:0] io_in_a_102,
  input  [31:0] io_in_a_103,
  input  [31:0] io_in_a_104,
  input  [31:0] io_in_a_105,
  input  [31:0] io_in_a_106,
  input  [31:0] io_in_a_107,
  input  [31:0] io_in_a_108,
  input  [31:0] io_in_a_109,
  input  [31:0] io_in_a_110,
  input  [31:0] io_in_a_111,
  input  [31:0] io_in_a_112,
  input  [31:0] io_in_a_113,
  input  [31:0] io_in_a_114,
  input  [31:0] io_in_a_115,
  input  [31:0] io_in_a_116,
  input  [31:0] io_in_a_117,
  input  [31:0] io_in_a_118,
  input  [31:0] io_in_a_119,
  input  [31:0] io_in_a_120,
  input  [31:0] io_in_a_121,
  input  [31:0] io_in_a_122,
  input  [31:0] io_in_a_123,
  input  [31:0] io_in_a_124,
  input  [31:0] io_in_a_125,
  input  [31:0] io_in_a_126,
  input  [31:0] io_in_a_127,
  input  [31:0] io_in_b_0,
  input  [31:0] io_in_b_1,
  input  [31:0] io_in_b_2,
  input  [31:0] io_in_b_3,
  input  [31:0] io_in_b_4,
  input  [31:0] io_in_b_5,
  input  [31:0] io_in_b_6,
  input  [31:0] io_in_b_7,
  input  [31:0] io_in_b_8,
  input  [31:0] io_in_b_9,
  input  [31:0] io_in_b_10,
  input  [31:0] io_in_b_11,
  input  [31:0] io_in_b_12,
  input  [31:0] io_in_b_13,
  input  [31:0] io_in_b_14,
  input  [31:0] io_in_b_15,
  input  [31:0] io_in_b_16,
  input  [31:0] io_in_b_17,
  input  [31:0] io_in_b_18,
  input  [31:0] io_in_b_19,
  input  [31:0] io_in_b_20,
  input  [31:0] io_in_b_21,
  input  [31:0] io_in_b_22,
  input  [31:0] io_in_b_23,
  input  [31:0] io_in_b_24,
  input  [31:0] io_in_b_25,
  input  [31:0] io_in_b_26,
  input  [31:0] io_in_b_27,
  input  [31:0] io_in_b_28,
  input  [31:0] io_in_b_29,
  input  [31:0] io_in_b_30,
  input  [31:0] io_in_b_31,
  input  [31:0] io_in_b_32,
  input  [31:0] io_in_b_33,
  input  [31:0] io_in_b_34,
  input  [31:0] io_in_b_35,
  input  [31:0] io_in_b_36,
  input  [31:0] io_in_b_37,
  input  [31:0] io_in_b_38,
  input  [31:0] io_in_b_39,
  input  [31:0] io_in_b_40,
  input  [31:0] io_in_b_41,
  input  [31:0] io_in_b_42,
  input  [31:0] io_in_b_43,
  input  [31:0] io_in_b_44,
  input  [31:0] io_in_b_45,
  input  [31:0] io_in_b_46,
  input  [31:0] io_in_b_47,
  input  [31:0] io_in_b_48,
  input  [31:0] io_in_b_49,
  input  [31:0] io_in_b_50,
  input  [31:0] io_in_b_51,
  input  [31:0] io_in_b_52,
  input  [31:0] io_in_b_53,
  input  [31:0] io_in_b_54,
  input  [31:0] io_in_b_55,
  input  [31:0] io_in_b_56,
  input  [31:0] io_in_b_57,
  input  [31:0] io_in_b_58,
  input  [31:0] io_in_b_59,
  input  [31:0] io_in_b_60,
  input  [31:0] io_in_b_61,
  input  [31:0] io_in_b_62,
  input  [31:0] io_in_b_63,
  input  [31:0] io_in_b_64,
  input  [31:0] io_in_b_65,
  input  [31:0] io_in_b_66,
  input  [31:0] io_in_b_67,
  input  [31:0] io_in_b_68,
  input  [31:0] io_in_b_69,
  input  [31:0] io_in_b_70,
  input  [31:0] io_in_b_71,
  input  [31:0] io_in_b_72,
  input  [31:0] io_in_b_73,
  input  [31:0] io_in_b_74,
  input  [31:0] io_in_b_75,
  input  [31:0] io_in_b_76,
  input  [31:0] io_in_b_77,
  input  [31:0] io_in_b_78,
  input  [31:0] io_in_b_79,
  input  [31:0] io_in_b_80,
  input  [31:0] io_in_b_81,
  input  [31:0] io_in_b_82,
  input  [31:0] io_in_b_83,
  input  [31:0] io_in_b_84,
  input  [31:0] io_in_b_85,
  input  [31:0] io_in_b_86,
  input  [31:0] io_in_b_87,
  input  [31:0] io_in_b_88,
  input  [31:0] io_in_b_89,
  input  [31:0] io_in_b_90,
  input  [31:0] io_in_b_91,
  input  [31:0] io_in_b_92,
  input  [31:0] io_in_b_93,
  input  [31:0] io_in_b_94,
  input  [31:0] io_in_b_95,
  input  [31:0] io_in_b_96,
  input  [31:0] io_in_b_97,
  input  [31:0] io_in_b_98,
  input  [31:0] io_in_b_99,
  input  [31:0] io_in_b_100,
  input  [31:0] io_in_b_101,
  input  [31:0] io_in_b_102,
  input  [31:0] io_in_b_103,
  input  [31:0] io_in_b_104,
  input  [31:0] io_in_b_105,
  input  [31:0] io_in_b_106,
  input  [31:0] io_in_b_107,
  input  [31:0] io_in_b_108,
  input  [31:0] io_in_b_109,
  input  [31:0] io_in_b_110,
  input  [31:0] io_in_b_111,
  input  [31:0] io_in_b_112,
  input  [31:0] io_in_b_113,
  input  [31:0] io_in_b_114,
  input  [31:0] io_in_b_115,
  input  [31:0] io_in_b_116,
  input  [31:0] io_in_b_117,
  input  [31:0] io_in_b_118,
  input  [31:0] io_in_b_119,
  input  [31:0] io_in_b_120,
  input  [31:0] io_in_b_121,
  input  [31:0] io_in_b_122,
  input  [31:0] io_in_b_123,
  input  [31:0] io_in_b_124,
  input  [31:0] io_in_b_125,
  input  [31:0] io_in_b_126,
  input  [31:0] io_in_b_127,
  output [31:0] io_out_s
);
  wire  FP_multiplier_10ccs_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_1_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_1_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_1_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_1_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_2_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_2_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_2_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_2_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_3_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_3_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_3_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_3_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_4_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_4_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_4_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_4_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_5_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_5_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_5_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_5_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_6_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_6_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_6_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_6_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_7_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_7_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_7_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_7_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_8_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_8_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_8_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_8_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_9_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_9_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_9_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_9_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_10_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_10_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_10_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_10_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_11_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_11_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_11_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_11_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_12_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_12_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_12_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_12_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_13_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_13_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_13_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_13_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_14_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_14_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_14_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_14_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_15_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_15_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_15_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_15_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_16_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_16_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_16_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_16_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_17_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_17_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_17_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_17_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_18_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_18_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_18_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_18_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_19_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_19_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_19_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_19_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_20_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_20_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_20_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_20_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_21_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_21_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_21_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_21_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_22_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_22_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_22_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_22_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_23_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_23_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_23_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_23_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_24_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_24_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_24_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_24_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_25_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_25_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_25_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_25_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_26_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_26_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_26_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_26_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_27_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_27_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_27_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_27_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_28_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_28_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_28_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_28_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_29_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_29_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_29_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_29_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_30_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_30_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_30_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_30_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_31_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_31_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_31_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_31_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_32_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_32_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_32_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_32_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_33_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_33_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_33_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_33_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_34_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_34_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_34_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_34_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_35_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_35_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_35_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_35_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_36_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_36_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_36_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_36_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_37_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_37_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_37_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_37_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_38_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_38_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_38_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_38_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_39_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_39_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_39_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_39_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_40_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_40_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_40_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_40_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_41_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_41_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_41_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_41_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_42_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_42_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_42_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_42_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_43_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_43_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_43_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_43_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_44_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_44_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_44_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_44_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_45_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_45_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_45_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_45_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_46_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_46_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_46_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_46_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_47_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_47_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_47_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_47_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_47_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_48_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_48_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_48_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_48_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_49_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_49_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_49_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_49_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_50_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_50_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_50_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_50_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_51_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_51_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_51_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_51_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_52_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_52_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_52_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_52_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_53_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_53_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_53_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_53_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_54_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_54_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_54_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_54_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_55_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_55_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_55_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_55_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_56_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_56_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_56_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_56_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_57_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_57_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_57_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_57_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_58_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_58_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_58_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_58_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_59_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_59_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_59_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_59_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_60_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_60_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_60_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_60_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_61_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_61_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_61_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_61_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_62_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_62_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_62_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_62_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_63_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_63_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_63_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_63_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_63_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_64_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_64_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_64_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_64_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_64_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_65_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_65_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_65_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_65_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_65_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_66_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_66_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_66_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_66_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_66_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_67_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_67_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_67_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_67_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_67_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_68_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_68_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_68_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_68_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_68_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_69_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_69_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_69_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_69_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_69_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_70_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_70_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_70_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_70_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_70_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_71_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_71_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_71_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_71_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_71_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_72_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_72_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_72_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_72_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_72_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_73_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_73_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_73_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_73_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_73_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_74_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_74_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_74_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_74_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_74_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_75_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_75_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_75_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_75_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_75_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_76_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_76_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_76_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_76_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_76_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_77_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_77_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_77_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_77_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_77_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_78_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_78_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_78_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_78_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_78_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_79_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_79_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_79_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_79_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_79_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_80_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_80_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_80_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_80_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_80_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_81_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_81_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_81_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_81_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_81_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_82_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_82_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_82_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_82_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_82_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_83_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_83_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_83_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_83_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_83_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_84_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_84_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_84_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_84_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_84_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_85_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_85_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_85_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_85_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_85_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_86_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_86_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_86_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_86_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_86_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_87_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_87_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_87_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_87_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_87_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_88_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_88_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_88_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_88_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_88_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_89_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_89_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_89_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_89_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_89_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_90_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_90_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_90_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_90_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_90_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_91_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_91_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_91_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_91_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_91_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_92_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_92_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_92_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_92_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_92_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_93_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_93_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_93_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_93_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_93_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_94_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_94_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_94_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_94_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_94_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_95_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_95_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_95_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_95_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_95_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_96_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_96_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_96_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_96_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_96_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_97_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_97_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_97_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_97_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_97_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_98_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_98_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_98_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_98_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_98_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_99_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_99_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_99_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_99_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_99_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_100_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_100_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_100_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_100_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_100_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_101_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_101_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_101_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_101_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_101_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_102_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_102_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_102_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_102_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_102_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_103_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_103_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_103_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_103_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_103_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_104_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_104_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_104_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_104_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_104_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_105_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_105_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_105_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_105_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_105_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_106_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_106_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_106_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_106_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_106_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_107_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_107_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_107_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_107_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_107_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_108_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_108_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_108_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_108_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_108_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_109_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_109_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_109_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_109_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_109_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_110_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_110_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_110_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_110_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_110_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_111_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_111_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_111_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_111_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_111_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_112_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_112_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_112_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_112_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_112_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_113_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_113_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_113_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_113_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_113_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_114_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_114_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_114_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_114_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_114_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_115_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_115_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_115_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_115_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_115_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_116_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_116_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_116_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_116_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_116_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_117_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_117_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_117_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_117_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_117_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_118_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_118_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_118_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_118_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_118_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_119_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_119_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_119_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_119_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_119_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_120_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_120_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_120_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_120_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_120_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_121_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_121_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_121_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_121_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_121_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_122_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_122_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_122_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_122_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_122_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_123_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_123_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_123_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_123_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_123_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_124_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_124_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_124_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_124_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_124_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_125_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_125_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_125_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_125_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_125_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_126_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_126_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_126_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_126_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_126_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_127_clock; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_multiplier_10ccs_127_reset; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_127_io_in_a; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_127_io_in_b; // @[FloatingPointDesigns.scala 2409:44]
  wire [31:0] FP_multiplier_10ccs_127_io_out_s; // @[FloatingPointDesigns.scala 2409:44]
  wire  FP_adder_13ccs_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_1_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_1_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_1_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_1_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_2_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_2_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_2_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_2_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_3_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_3_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_3_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_3_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_4_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_4_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_4_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_4_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_5_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_5_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_5_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_5_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_6_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_6_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_6_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_6_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_7_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_7_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_7_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_7_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_8_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_8_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_8_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_8_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_9_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_9_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_9_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_9_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_10_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_10_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_10_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_10_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_11_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_11_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_11_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_11_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_12_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_12_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_12_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_12_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_13_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_13_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_13_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_13_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_14_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_14_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_14_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_14_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_15_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_15_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_15_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_15_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_16_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_16_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_16_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_16_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_17_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_17_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_17_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_17_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_18_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_18_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_18_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_18_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_19_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_19_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_19_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_19_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_20_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_20_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_20_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_20_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_21_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_21_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_21_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_21_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_22_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_22_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_22_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_22_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_23_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_23_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_23_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_23_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_24_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_24_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_24_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_24_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_25_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_25_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_25_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_25_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_26_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_26_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_26_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_26_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_27_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_27_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_27_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_27_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_28_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_28_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_28_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_28_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_29_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_29_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_29_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_29_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_30_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_30_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_30_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_30_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_31_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_31_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_31_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_31_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_32_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_32_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_32_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_32_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_33_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_33_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_33_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_33_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_34_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_34_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_34_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_34_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_35_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_35_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_35_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_35_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_36_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_36_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_36_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_36_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_37_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_37_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_37_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_37_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_38_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_38_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_38_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_38_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_39_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_39_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_39_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_39_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_40_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_40_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_40_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_40_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_41_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_41_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_41_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_41_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_42_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_42_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_42_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_42_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_43_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_43_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_43_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_43_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_44_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_44_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_44_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_44_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_45_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_45_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_45_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_45_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_46_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_46_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_46_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_46_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_47_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_47_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_47_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_47_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_47_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_48_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_48_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_48_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_48_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_49_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_49_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_49_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_49_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_50_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_50_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_50_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_50_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_51_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_51_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_51_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_51_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_52_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_52_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_52_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_52_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_53_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_53_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_53_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_53_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_54_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_54_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_54_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_54_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_55_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_55_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_55_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_55_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_56_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_56_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_56_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_56_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_57_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_57_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_57_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_57_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_58_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_58_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_58_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_58_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_59_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_59_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_59_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_59_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_60_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_60_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_60_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_60_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_61_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_61_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_61_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_61_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_62_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_62_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_62_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_62_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_63_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_63_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_63_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_63_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_63_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_64_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_64_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_64_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_64_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_64_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_65_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_65_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_65_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_65_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_65_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_66_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_66_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_66_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_66_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_66_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_67_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_67_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_67_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_67_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_67_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_68_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_68_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_68_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_68_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_68_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_69_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_69_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_69_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_69_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_69_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_70_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_70_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_70_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_70_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_70_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_71_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_71_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_71_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_71_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_71_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_72_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_72_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_72_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_72_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_72_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_73_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_73_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_73_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_73_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_73_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_74_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_74_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_74_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_74_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_74_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_75_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_75_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_75_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_75_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_75_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_76_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_76_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_76_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_76_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_76_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_77_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_77_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_77_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_77_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_77_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_78_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_78_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_78_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_78_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_78_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_79_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_79_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_79_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_79_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_79_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_80_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_80_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_80_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_80_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_80_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_81_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_81_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_81_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_81_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_81_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_82_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_82_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_82_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_82_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_82_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_83_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_83_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_83_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_83_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_83_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_84_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_84_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_84_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_84_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_84_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_85_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_85_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_85_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_85_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_85_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_86_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_86_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_86_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_86_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_86_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_87_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_87_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_87_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_87_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_87_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_88_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_88_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_88_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_88_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_88_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_89_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_89_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_89_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_89_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_89_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_90_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_90_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_90_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_90_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_90_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_91_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_91_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_91_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_91_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_91_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_92_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_92_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_92_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_92_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_92_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_93_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_93_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_93_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_93_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_93_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_94_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_94_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_94_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_94_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_94_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_95_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_95_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_95_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_95_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_95_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_96_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_96_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_96_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_96_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_96_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_97_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_97_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_97_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_97_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_97_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_98_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_98_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_98_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_98_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_98_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_99_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_99_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_99_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_99_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_99_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_100_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_100_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_100_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_100_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_100_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_101_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_101_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_101_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_101_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_101_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_102_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_102_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_102_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_102_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_102_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_103_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_103_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_103_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_103_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_103_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_104_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_104_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_104_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_104_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_104_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_105_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_105_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_105_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_105_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_105_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_106_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_106_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_106_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_106_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_106_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_107_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_107_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_107_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_107_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_107_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_108_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_108_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_108_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_108_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_108_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_109_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_109_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_109_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_109_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_109_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_110_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_110_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_110_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_110_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_110_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_111_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_111_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_111_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_111_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_111_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_112_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_112_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_112_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_112_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_112_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_113_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_113_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_113_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_113_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_113_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_114_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_114_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_114_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_114_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_114_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_115_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_115_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_115_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_115_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_115_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_116_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_116_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_116_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_116_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_116_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_117_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_117_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_117_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_117_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_117_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_118_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_118_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_118_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_118_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_118_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_119_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_119_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_119_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_119_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_119_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_120_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_120_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_120_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_120_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_120_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_121_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_121_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_121_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_121_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_121_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_122_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_122_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_122_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_122_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_122_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_123_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_123_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_123_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_123_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_123_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_124_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_124_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_124_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_124_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_124_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_125_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_125_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_125_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_125_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_125_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_126_clock; // @[FloatingPointDesigns.scala 2417:17]
  wire  FP_adder_13ccs_126_reset; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_126_io_in_a; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_126_io_in_b; // @[FloatingPointDesigns.scala 2417:17]
  wire [31:0] FP_adder_13ccs_126_io_out_s; // @[FloatingPointDesigns.scala 2417:17]
  FP_multiplier_10ccs FP_multiplier_10ccs ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_clock),
    .reset(FP_multiplier_10ccs_reset),
    .io_in_a(FP_multiplier_10ccs_io_in_a),
    .io_in_b(FP_multiplier_10ccs_io_in_b),
    .io_out_s(FP_multiplier_10ccs_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_1 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_1_clock),
    .reset(FP_multiplier_10ccs_1_reset),
    .io_in_a(FP_multiplier_10ccs_1_io_in_a),
    .io_in_b(FP_multiplier_10ccs_1_io_in_b),
    .io_out_s(FP_multiplier_10ccs_1_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_2 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_2_clock),
    .reset(FP_multiplier_10ccs_2_reset),
    .io_in_a(FP_multiplier_10ccs_2_io_in_a),
    .io_in_b(FP_multiplier_10ccs_2_io_in_b),
    .io_out_s(FP_multiplier_10ccs_2_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_3 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_3_clock),
    .reset(FP_multiplier_10ccs_3_reset),
    .io_in_a(FP_multiplier_10ccs_3_io_in_a),
    .io_in_b(FP_multiplier_10ccs_3_io_in_b),
    .io_out_s(FP_multiplier_10ccs_3_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_4 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_4_clock),
    .reset(FP_multiplier_10ccs_4_reset),
    .io_in_a(FP_multiplier_10ccs_4_io_in_a),
    .io_in_b(FP_multiplier_10ccs_4_io_in_b),
    .io_out_s(FP_multiplier_10ccs_4_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_5 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_5_clock),
    .reset(FP_multiplier_10ccs_5_reset),
    .io_in_a(FP_multiplier_10ccs_5_io_in_a),
    .io_in_b(FP_multiplier_10ccs_5_io_in_b),
    .io_out_s(FP_multiplier_10ccs_5_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_6 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_6_clock),
    .reset(FP_multiplier_10ccs_6_reset),
    .io_in_a(FP_multiplier_10ccs_6_io_in_a),
    .io_in_b(FP_multiplier_10ccs_6_io_in_b),
    .io_out_s(FP_multiplier_10ccs_6_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_7 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_7_clock),
    .reset(FP_multiplier_10ccs_7_reset),
    .io_in_a(FP_multiplier_10ccs_7_io_in_a),
    .io_in_b(FP_multiplier_10ccs_7_io_in_b),
    .io_out_s(FP_multiplier_10ccs_7_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_8 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_8_clock),
    .reset(FP_multiplier_10ccs_8_reset),
    .io_in_a(FP_multiplier_10ccs_8_io_in_a),
    .io_in_b(FP_multiplier_10ccs_8_io_in_b),
    .io_out_s(FP_multiplier_10ccs_8_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_9 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_9_clock),
    .reset(FP_multiplier_10ccs_9_reset),
    .io_in_a(FP_multiplier_10ccs_9_io_in_a),
    .io_in_b(FP_multiplier_10ccs_9_io_in_b),
    .io_out_s(FP_multiplier_10ccs_9_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_10 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_10_clock),
    .reset(FP_multiplier_10ccs_10_reset),
    .io_in_a(FP_multiplier_10ccs_10_io_in_a),
    .io_in_b(FP_multiplier_10ccs_10_io_in_b),
    .io_out_s(FP_multiplier_10ccs_10_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_11 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_11_clock),
    .reset(FP_multiplier_10ccs_11_reset),
    .io_in_a(FP_multiplier_10ccs_11_io_in_a),
    .io_in_b(FP_multiplier_10ccs_11_io_in_b),
    .io_out_s(FP_multiplier_10ccs_11_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_12 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_12_clock),
    .reset(FP_multiplier_10ccs_12_reset),
    .io_in_a(FP_multiplier_10ccs_12_io_in_a),
    .io_in_b(FP_multiplier_10ccs_12_io_in_b),
    .io_out_s(FP_multiplier_10ccs_12_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_13 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_13_clock),
    .reset(FP_multiplier_10ccs_13_reset),
    .io_in_a(FP_multiplier_10ccs_13_io_in_a),
    .io_in_b(FP_multiplier_10ccs_13_io_in_b),
    .io_out_s(FP_multiplier_10ccs_13_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_14 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_14_clock),
    .reset(FP_multiplier_10ccs_14_reset),
    .io_in_a(FP_multiplier_10ccs_14_io_in_a),
    .io_in_b(FP_multiplier_10ccs_14_io_in_b),
    .io_out_s(FP_multiplier_10ccs_14_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_15 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_15_clock),
    .reset(FP_multiplier_10ccs_15_reset),
    .io_in_a(FP_multiplier_10ccs_15_io_in_a),
    .io_in_b(FP_multiplier_10ccs_15_io_in_b),
    .io_out_s(FP_multiplier_10ccs_15_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_16 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_16_clock),
    .reset(FP_multiplier_10ccs_16_reset),
    .io_in_a(FP_multiplier_10ccs_16_io_in_a),
    .io_in_b(FP_multiplier_10ccs_16_io_in_b),
    .io_out_s(FP_multiplier_10ccs_16_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_17 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_17_clock),
    .reset(FP_multiplier_10ccs_17_reset),
    .io_in_a(FP_multiplier_10ccs_17_io_in_a),
    .io_in_b(FP_multiplier_10ccs_17_io_in_b),
    .io_out_s(FP_multiplier_10ccs_17_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_18 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_18_clock),
    .reset(FP_multiplier_10ccs_18_reset),
    .io_in_a(FP_multiplier_10ccs_18_io_in_a),
    .io_in_b(FP_multiplier_10ccs_18_io_in_b),
    .io_out_s(FP_multiplier_10ccs_18_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_19 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_19_clock),
    .reset(FP_multiplier_10ccs_19_reset),
    .io_in_a(FP_multiplier_10ccs_19_io_in_a),
    .io_in_b(FP_multiplier_10ccs_19_io_in_b),
    .io_out_s(FP_multiplier_10ccs_19_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_20 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_20_clock),
    .reset(FP_multiplier_10ccs_20_reset),
    .io_in_a(FP_multiplier_10ccs_20_io_in_a),
    .io_in_b(FP_multiplier_10ccs_20_io_in_b),
    .io_out_s(FP_multiplier_10ccs_20_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_21 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_21_clock),
    .reset(FP_multiplier_10ccs_21_reset),
    .io_in_a(FP_multiplier_10ccs_21_io_in_a),
    .io_in_b(FP_multiplier_10ccs_21_io_in_b),
    .io_out_s(FP_multiplier_10ccs_21_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_22 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_22_clock),
    .reset(FP_multiplier_10ccs_22_reset),
    .io_in_a(FP_multiplier_10ccs_22_io_in_a),
    .io_in_b(FP_multiplier_10ccs_22_io_in_b),
    .io_out_s(FP_multiplier_10ccs_22_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_23 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_23_clock),
    .reset(FP_multiplier_10ccs_23_reset),
    .io_in_a(FP_multiplier_10ccs_23_io_in_a),
    .io_in_b(FP_multiplier_10ccs_23_io_in_b),
    .io_out_s(FP_multiplier_10ccs_23_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_24 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_24_clock),
    .reset(FP_multiplier_10ccs_24_reset),
    .io_in_a(FP_multiplier_10ccs_24_io_in_a),
    .io_in_b(FP_multiplier_10ccs_24_io_in_b),
    .io_out_s(FP_multiplier_10ccs_24_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_25 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_25_clock),
    .reset(FP_multiplier_10ccs_25_reset),
    .io_in_a(FP_multiplier_10ccs_25_io_in_a),
    .io_in_b(FP_multiplier_10ccs_25_io_in_b),
    .io_out_s(FP_multiplier_10ccs_25_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_26 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_26_clock),
    .reset(FP_multiplier_10ccs_26_reset),
    .io_in_a(FP_multiplier_10ccs_26_io_in_a),
    .io_in_b(FP_multiplier_10ccs_26_io_in_b),
    .io_out_s(FP_multiplier_10ccs_26_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_27 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_27_clock),
    .reset(FP_multiplier_10ccs_27_reset),
    .io_in_a(FP_multiplier_10ccs_27_io_in_a),
    .io_in_b(FP_multiplier_10ccs_27_io_in_b),
    .io_out_s(FP_multiplier_10ccs_27_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_28 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_28_clock),
    .reset(FP_multiplier_10ccs_28_reset),
    .io_in_a(FP_multiplier_10ccs_28_io_in_a),
    .io_in_b(FP_multiplier_10ccs_28_io_in_b),
    .io_out_s(FP_multiplier_10ccs_28_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_29 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_29_clock),
    .reset(FP_multiplier_10ccs_29_reset),
    .io_in_a(FP_multiplier_10ccs_29_io_in_a),
    .io_in_b(FP_multiplier_10ccs_29_io_in_b),
    .io_out_s(FP_multiplier_10ccs_29_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_30 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_30_clock),
    .reset(FP_multiplier_10ccs_30_reset),
    .io_in_a(FP_multiplier_10ccs_30_io_in_a),
    .io_in_b(FP_multiplier_10ccs_30_io_in_b),
    .io_out_s(FP_multiplier_10ccs_30_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_31 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_31_clock),
    .reset(FP_multiplier_10ccs_31_reset),
    .io_in_a(FP_multiplier_10ccs_31_io_in_a),
    .io_in_b(FP_multiplier_10ccs_31_io_in_b),
    .io_out_s(FP_multiplier_10ccs_31_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_32 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_32_clock),
    .reset(FP_multiplier_10ccs_32_reset),
    .io_in_a(FP_multiplier_10ccs_32_io_in_a),
    .io_in_b(FP_multiplier_10ccs_32_io_in_b),
    .io_out_s(FP_multiplier_10ccs_32_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_33 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_33_clock),
    .reset(FP_multiplier_10ccs_33_reset),
    .io_in_a(FP_multiplier_10ccs_33_io_in_a),
    .io_in_b(FP_multiplier_10ccs_33_io_in_b),
    .io_out_s(FP_multiplier_10ccs_33_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_34 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_34_clock),
    .reset(FP_multiplier_10ccs_34_reset),
    .io_in_a(FP_multiplier_10ccs_34_io_in_a),
    .io_in_b(FP_multiplier_10ccs_34_io_in_b),
    .io_out_s(FP_multiplier_10ccs_34_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_35 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_35_clock),
    .reset(FP_multiplier_10ccs_35_reset),
    .io_in_a(FP_multiplier_10ccs_35_io_in_a),
    .io_in_b(FP_multiplier_10ccs_35_io_in_b),
    .io_out_s(FP_multiplier_10ccs_35_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_36 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_36_clock),
    .reset(FP_multiplier_10ccs_36_reset),
    .io_in_a(FP_multiplier_10ccs_36_io_in_a),
    .io_in_b(FP_multiplier_10ccs_36_io_in_b),
    .io_out_s(FP_multiplier_10ccs_36_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_37 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_37_clock),
    .reset(FP_multiplier_10ccs_37_reset),
    .io_in_a(FP_multiplier_10ccs_37_io_in_a),
    .io_in_b(FP_multiplier_10ccs_37_io_in_b),
    .io_out_s(FP_multiplier_10ccs_37_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_38 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_38_clock),
    .reset(FP_multiplier_10ccs_38_reset),
    .io_in_a(FP_multiplier_10ccs_38_io_in_a),
    .io_in_b(FP_multiplier_10ccs_38_io_in_b),
    .io_out_s(FP_multiplier_10ccs_38_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_39 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_39_clock),
    .reset(FP_multiplier_10ccs_39_reset),
    .io_in_a(FP_multiplier_10ccs_39_io_in_a),
    .io_in_b(FP_multiplier_10ccs_39_io_in_b),
    .io_out_s(FP_multiplier_10ccs_39_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_40 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_40_clock),
    .reset(FP_multiplier_10ccs_40_reset),
    .io_in_a(FP_multiplier_10ccs_40_io_in_a),
    .io_in_b(FP_multiplier_10ccs_40_io_in_b),
    .io_out_s(FP_multiplier_10ccs_40_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_41 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_41_clock),
    .reset(FP_multiplier_10ccs_41_reset),
    .io_in_a(FP_multiplier_10ccs_41_io_in_a),
    .io_in_b(FP_multiplier_10ccs_41_io_in_b),
    .io_out_s(FP_multiplier_10ccs_41_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_42 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_42_clock),
    .reset(FP_multiplier_10ccs_42_reset),
    .io_in_a(FP_multiplier_10ccs_42_io_in_a),
    .io_in_b(FP_multiplier_10ccs_42_io_in_b),
    .io_out_s(FP_multiplier_10ccs_42_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_43 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_43_clock),
    .reset(FP_multiplier_10ccs_43_reset),
    .io_in_a(FP_multiplier_10ccs_43_io_in_a),
    .io_in_b(FP_multiplier_10ccs_43_io_in_b),
    .io_out_s(FP_multiplier_10ccs_43_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_44 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_44_clock),
    .reset(FP_multiplier_10ccs_44_reset),
    .io_in_a(FP_multiplier_10ccs_44_io_in_a),
    .io_in_b(FP_multiplier_10ccs_44_io_in_b),
    .io_out_s(FP_multiplier_10ccs_44_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_45 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_45_clock),
    .reset(FP_multiplier_10ccs_45_reset),
    .io_in_a(FP_multiplier_10ccs_45_io_in_a),
    .io_in_b(FP_multiplier_10ccs_45_io_in_b),
    .io_out_s(FP_multiplier_10ccs_45_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_46 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_46_clock),
    .reset(FP_multiplier_10ccs_46_reset),
    .io_in_a(FP_multiplier_10ccs_46_io_in_a),
    .io_in_b(FP_multiplier_10ccs_46_io_in_b),
    .io_out_s(FP_multiplier_10ccs_46_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_47 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_47_clock),
    .reset(FP_multiplier_10ccs_47_reset),
    .io_in_a(FP_multiplier_10ccs_47_io_in_a),
    .io_in_b(FP_multiplier_10ccs_47_io_in_b),
    .io_out_s(FP_multiplier_10ccs_47_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_48 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_48_clock),
    .reset(FP_multiplier_10ccs_48_reset),
    .io_in_a(FP_multiplier_10ccs_48_io_in_a),
    .io_in_b(FP_multiplier_10ccs_48_io_in_b),
    .io_out_s(FP_multiplier_10ccs_48_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_49 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_49_clock),
    .reset(FP_multiplier_10ccs_49_reset),
    .io_in_a(FP_multiplier_10ccs_49_io_in_a),
    .io_in_b(FP_multiplier_10ccs_49_io_in_b),
    .io_out_s(FP_multiplier_10ccs_49_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_50 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_50_clock),
    .reset(FP_multiplier_10ccs_50_reset),
    .io_in_a(FP_multiplier_10ccs_50_io_in_a),
    .io_in_b(FP_multiplier_10ccs_50_io_in_b),
    .io_out_s(FP_multiplier_10ccs_50_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_51 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_51_clock),
    .reset(FP_multiplier_10ccs_51_reset),
    .io_in_a(FP_multiplier_10ccs_51_io_in_a),
    .io_in_b(FP_multiplier_10ccs_51_io_in_b),
    .io_out_s(FP_multiplier_10ccs_51_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_52 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_52_clock),
    .reset(FP_multiplier_10ccs_52_reset),
    .io_in_a(FP_multiplier_10ccs_52_io_in_a),
    .io_in_b(FP_multiplier_10ccs_52_io_in_b),
    .io_out_s(FP_multiplier_10ccs_52_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_53 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_53_clock),
    .reset(FP_multiplier_10ccs_53_reset),
    .io_in_a(FP_multiplier_10ccs_53_io_in_a),
    .io_in_b(FP_multiplier_10ccs_53_io_in_b),
    .io_out_s(FP_multiplier_10ccs_53_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_54 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_54_clock),
    .reset(FP_multiplier_10ccs_54_reset),
    .io_in_a(FP_multiplier_10ccs_54_io_in_a),
    .io_in_b(FP_multiplier_10ccs_54_io_in_b),
    .io_out_s(FP_multiplier_10ccs_54_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_55 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_55_clock),
    .reset(FP_multiplier_10ccs_55_reset),
    .io_in_a(FP_multiplier_10ccs_55_io_in_a),
    .io_in_b(FP_multiplier_10ccs_55_io_in_b),
    .io_out_s(FP_multiplier_10ccs_55_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_56 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_56_clock),
    .reset(FP_multiplier_10ccs_56_reset),
    .io_in_a(FP_multiplier_10ccs_56_io_in_a),
    .io_in_b(FP_multiplier_10ccs_56_io_in_b),
    .io_out_s(FP_multiplier_10ccs_56_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_57 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_57_clock),
    .reset(FP_multiplier_10ccs_57_reset),
    .io_in_a(FP_multiplier_10ccs_57_io_in_a),
    .io_in_b(FP_multiplier_10ccs_57_io_in_b),
    .io_out_s(FP_multiplier_10ccs_57_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_58 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_58_clock),
    .reset(FP_multiplier_10ccs_58_reset),
    .io_in_a(FP_multiplier_10ccs_58_io_in_a),
    .io_in_b(FP_multiplier_10ccs_58_io_in_b),
    .io_out_s(FP_multiplier_10ccs_58_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_59 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_59_clock),
    .reset(FP_multiplier_10ccs_59_reset),
    .io_in_a(FP_multiplier_10ccs_59_io_in_a),
    .io_in_b(FP_multiplier_10ccs_59_io_in_b),
    .io_out_s(FP_multiplier_10ccs_59_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_60 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_60_clock),
    .reset(FP_multiplier_10ccs_60_reset),
    .io_in_a(FP_multiplier_10ccs_60_io_in_a),
    .io_in_b(FP_multiplier_10ccs_60_io_in_b),
    .io_out_s(FP_multiplier_10ccs_60_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_61 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_61_clock),
    .reset(FP_multiplier_10ccs_61_reset),
    .io_in_a(FP_multiplier_10ccs_61_io_in_a),
    .io_in_b(FP_multiplier_10ccs_61_io_in_b),
    .io_out_s(FP_multiplier_10ccs_61_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_62 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_62_clock),
    .reset(FP_multiplier_10ccs_62_reset),
    .io_in_a(FP_multiplier_10ccs_62_io_in_a),
    .io_in_b(FP_multiplier_10ccs_62_io_in_b),
    .io_out_s(FP_multiplier_10ccs_62_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_63 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_63_clock),
    .reset(FP_multiplier_10ccs_63_reset),
    .io_in_a(FP_multiplier_10ccs_63_io_in_a),
    .io_in_b(FP_multiplier_10ccs_63_io_in_b),
    .io_out_s(FP_multiplier_10ccs_63_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_64 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_64_clock),
    .reset(FP_multiplier_10ccs_64_reset),
    .io_in_a(FP_multiplier_10ccs_64_io_in_a),
    .io_in_b(FP_multiplier_10ccs_64_io_in_b),
    .io_out_s(FP_multiplier_10ccs_64_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_65 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_65_clock),
    .reset(FP_multiplier_10ccs_65_reset),
    .io_in_a(FP_multiplier_10ccs_65_io_in_a),
    .io_in_b(FP_multiplier_10ccs_65_io_in_b),
    .io_out_s(FP_multiplier_10ccs_65_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_66 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_66_clock),
    .reset(FP_multiplier_10ccs_66_reset),
    .io_in_a(FP_multiplier_10ccs_66_io_in_a),
    .io_in_b(FP_multiplier_10ccs_66_io_in_b),
    .io_out_s(FP_multiplier_10ccs_66_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_67 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_67_clock),
    .reset(FP_multiplier_10ccs_67_reset),
    .io_in_a(FP_multiplier_10ccs_67_io_in_a),
    .io_in_b(FP_multiplier_10ccs_67_io_in_b),
    .io_out_s(FP_multiplier_10ccs_67_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_68 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_68_clock),
    .reset(FP_multiplier_10ccs_68_reset),
    .io_in_a(FP_multiplier_10ccs_68_io_in_a),
    .io_in_b(FP_multiplier_10ccs_68_io_in_b),
    .io_out_s(FP_multiplier_10ccs_68_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_69 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_69_clock),
    .reset(FP_multiplier_10ccs_69_reset),
    .io_in_a(FP_multiplier_10ccs_69_io_in_a),
    .io_in_b(FP_multiplier_10ccs_69_io_in_b),
    .io_out_s(FP_multiplier_10ccs_69_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_70 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_70_clock),
    .reset(FP_multiplier_10ccs_70_reset),
    .io_in_a(FP_multiplier_10ccs_70_io_in_a),
    .io_in_b(FP_multiplier_10ccs_70_io_in_b),
    .io_out_s(FP_multiplier_10ccs_70_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_71 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_71_clock),
    .reset(FP_multiplier_10ccs_71_reset),
    .io_in_a(FP_multiplier_10ccs_71_io_in_a),
    .io_in_b(FP_multiplier_10ccs_71_io_in_b),
    .io_out_s(FP_multiplier_10ccs_71_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_72 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_72_clock),
    .reset(FP_multiplier_10ccs_72_reset),
    .io_in_a(FP_multiplier_10ccs_72_io_in_a),
    .io_in_b(FP_multiplier_10ccs_72_io_in_b),
    .io_out_s(FP_multiplier_10ccs_72_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_73 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_73_clock),
    .reset(FP_multiplier_10ccs_73_reset),
    .io_in_a(FP_multiplier_10ccs_73_io_in_a),
    .io_in_b(FP_multiplier_10ccs_73_io_in_b),
    .io_out_s(FP_multiplier_10ccs_73_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_74 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_74_clock),
    .reset(FP_multiplier_10ccs_74_reset),
    .io_in_a(FP_multiplier_10ccs_74_io_in_a),
    .io_in_b(FP_multiplier_10ccs_74_io_in_b),
    .io_out_s(FP_multiplier_10ccs_74_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_75 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_75_clock),
    .reset(FP_multiplier_10ccs_75_reset),
    .io_in_a(FP_multiplier_10ccs_75_io_in_a),
    .io_in_b(FP_multiplier_10ccs_75_io_in_b),
    .io_out_s(FP_multiplier_10ccs_75_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_76 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_76_clock),
    .reset(FP_multiplier_10ccs_76_reset),
    .io_in_a(FP_multiplier_10ccs_76_io_in_a),
    .io_in_b(FP_multiplier_10ccs_76_io_in_b),
    .io_out_s(FP_multiplier_10ccs_76_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_77 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_77_clock),
    .reset(FP_multiplier_10ccs_77_reset),
    .io_in_a(FP_multiplier_10ccs_77_io_in_a),
    .io_in_b(FP_multiplier_10ccs_77_io_in_b),
    .io_out_s(FP_multiplier_10ccs_77_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_78 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_78_clock),
    .reset(FP_multiplier_10ccs_78_reset),
    .io_in_a(FP_multiplier_10ccs_78_io_in_a),
    .io_in_b(FP_multiplier_10ccs_78_io_in_b),
    .io_out_s(FP_multiplier_10ccs_78_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_79 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_79_clock),
    .reset(FP_multiplier_10ccs_79_reset),
    .io_in_a(FP_multiplier_10ccs_79_io_in_a),
    .io_in_b(FP_multiplier_10ccs_79_io_in_b),
    .io_out_s(FP_multiplier_10ccs_79_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_80 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_80_clock),
    .reset(FP_multiplier_10ccs_80_reset),
    .io_in_a(FP_multiplier_10ccs_80_io_in_a),
    .io_in_b(FP_multiplier_10ccs_80_io_in_b),
    .io_out_s(FP_multiplier_10ccs_80_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_81 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_81_clock),
    .reset(FP_multiplier_10ccs_81_reset),
    .io_in_a(FP_multiplier_10ccs_81_io_in_a),
    .io_in_b(FP_multiplier_10ccs_81_io_in_b),
    .io_out_s(FP_multiplier_10ccs_81_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_82 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_82_clock),
    .reset(FP_multiplier_10ccs_82_reset),
    .io_in_a(FP_multiplier_10ccs_82_io_in_a),
    .io_in_b(FP_multiplier_10ccs_82_io_in_b),
    .io_out_s(FP_multiplier_10ccs_82_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_83 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_83_clock),
    .reset(FP_multiplier_10ccs_83_reset),
    .io_in_a(FP_multiplier_10ccs_83_io_in_a),
    .io_in_b(FP_multiplier_10ccs_83_io_in_b),
    .io_out_s(FP_multiplier_10ccs_83_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_84 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_84_clock),
    .reset(FP_multiplier_10ccs_84_reset),
    .io_in_a(FP_multiplier_10ccs_84_io_in_a),
    .io_in_b(FP_multiplier_10ccs_84_io_in_b),
    .io_out_s(FP_multiplier_10ccs_84_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_85 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_85_clock),
    .reset(FP_multiplier_10ccs_85_reset),
    .io_in_a(FP_multiplier_10ccs_85_io_in_a),
    .io_in_b(FP_multiplier_10ccs_85_io_in_b),
    .io_out_s(FP_multiplier_10ccs_85_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_86 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_86_clock),
    .reset(FP_multiplier_10ccs_86_reset),
    .io_in_a(FP_multiplier_10ccs_86_io_in_a),
    .io_in_b(FP_multiplier_10ccs_86_io_in_b),
    .io_out_s(FP_multiplier_10ccs_86_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_87 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_87_clock),
    .reset(FP_multiplier_10ccs_87_reset),
    .io_in_a(FP_multiplier_10ccs_87_io_in_a),
    .io_in_b(FP_multiplier_10ccs_87_io_in_b),
    .io_out_s(FP_multiplier_10ccs_87_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_88 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_88_clock),
    .reset(FP_multiplier_10ccs_88_reset),
    .io_in_a(FP_multiplier_10ccs_88_io_in_a),
    .io_in_b(FP_multiplier_10ccs_88_io_in_b),
    .io_out_s(FP_multiplier_10ccs_88_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_89 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_89_clock),
    .reset(FP_multiplier_10ccs_89_reset),
    .io_in_a(FP_multiplier_10ccs_89_io_in_a),
    .io_in_b(FP_multiplier_10ccs_89_io_in_b),
    .io_out_s(FP_multiplier_10ccs_89_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_90 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_90_clock),
    .reset(FP_multiplier_10ccs_90_reset),
    .io_in_a(FP_multiplier_10ccs_90_io_in_a),
    .io_in_b(FP_multiplier_10ccs_90_io_in_b),
    .io_out_s(FP_multiplier_10ccs_90_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_91 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_91_clock),
    .reset(FP_multiplier_10ccs_91_reset),
    .io_in_a(FP_multiplier_10ccs_91_io_in_a),
    .io_in_b(FP_multiplier_10ccs_91_io_in_b),
    .io_out_s(FP_multiplier_10ccs_91_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_92 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_92_clock),
    .reset(FP_multiplier_10ccs_92_reset),
    .io_in_a(FP_multiplier_10ccs_92_io_in_a),
    .io_in_b(FP_multiplier_10ccs_92_io_in_b),
    .io_out_s(FP_multiplier_10ccs_92_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_93 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_93_clock),
    .reset(FP_multiplier_10ccs_93_reset),
    .io_in_a(FP_multiplier_10ccs_93_io_in_a),
    .io_in_b(FP_multiplier_10ccs_93_io_in_b),
    .io_out_s(FP_multiplier_10ccs_93_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_94 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_94_clock),
    .reset(FP_multiplier_10ccs_94_reset),
    .io_in_a(FP_multiplier_10ccs_94_io_in_a),
    .io_in_b(FP_multiplier_10ccs_94_io_in_b),
    .io_out_s(FP_multiplier_10ccs_94_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_95 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_95_clock),
    .reset(FP_multiplier_10ccs_95_reset),
    .io_in_a(FP_multiplier_10ccs_95_io_in_a),
    .io_in_b(FP_multiplier_10ccs_95_io_in_b),
    .io_out_s(FP_multiplier_10ccs_95_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_96 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_96_clock),
    .reset(FP_multiplier_10ccs_96_reset),
    .io_in_a(FP_multiplier_10ccs_96_io_in_a),
    .io_in_b(FP_multiplier_10ccs_96_io_in_b),
    .io_out_s(FP_multiplier_10ccs_96_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_97 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_97_clock),
    .reset(FP_multiplier_10ccs_97_reset),
    .io_in_a(FP_multiplier_10ccs_97_io_in_a),
    .io_in_b(FP_multiplier_10ccs_97_io_in_b),
    .io_out_s(FP_multiplier_10ccs_97_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_98 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_98_clock),
    .reset(FP_multiplier_10ccs_98_reset),
    .io_in_a(FP_multiplier_10ccs_98_io_in_a),
    .io_in_b(FP_multiplier_10ccs_98_io_in_b),
    .io_out_s(FP_multiplier_10ccs_98_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_99 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_99_clock),
    .reset(FP_multiplier_10ccs_99_reset),
    .io_in_a(FP_multiplier_10ccs_99_io_in_a),
    .io_in_b(FP_multiplier_10ccs_99_io_in_b),
    .io_out_s(FP_multiplier_10ccs_99_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_100 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_100_clock),
    .reset(FP_multiplier_10ccs_100_reset),
    .io_in_a(FP_multiplier_10ccs_100_io_in_a),
    .io_in_b(FP_multiplier_10ccs_100_io_in_b),
    .io_out_s(FP_multiplier_10ccs_100_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_101 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_101_clock),
    .reset(FP_multiplier_10ccs_101_reset),
    .io_in_a(FP_multiplier_10ccs_101_io_in_a),
    .io_in_b(FP_multiplier_10ccs_101_io_in_b),
    .io_out_s(FP_multiplier_10ccs_101_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_102 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_102_clock),
    .reset(FP_multiplier_10ccs_102_reset),
    .io_in_a(FP_multiplier_10ccs_102_io_in_a),
    .io_in_b(FP_multiplier_10ccs_102_io_in_b),
    .io_out_s(FP_multiplier_10ccs_102_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_103 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_103_clock),
    .reset(FP_multiplier_10ccs_103_reset),
    .io_in_a(FP_multiplier_10ccs_103_io_in_a),
    .io_in_b(FP_multiplier_10ccs_103_io_in_b),
    .io_out_s(FP_multiplier_10ccs_103_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_104 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_104_clock),
    .reset(FP_multiplier_10ccs_104_reset),
    .io_in_a(FP_multiplier_10ccs_104_io_in_a),
    .io_in_b(FP_multiplier_10ccs_104_io_in_b),
    .io_out_s(FP_multiplier_10ccs_104_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_105 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_105_clock),
    .reset(FP_multiplier_10ccs_105_reset),
    .io_in_a(FP_multiplier_10ccs_105_io_in_a),
    .io_in_b(FP_multiplier_10ccs_105_io_in_b),
    .io_out_s(FP_multiplier_10ccs_105_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_106 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_106_clock),
    .reset(FP_multiplier_10ccs_106_reset),
    .io_in_a(FP_multiplier_10ccs_106_io_in_a),
    .io_in_b(FP_multiplier_10ccs_106_io_in_b),
    .io_out_s(FP_multiplier_10ccs_106_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_107 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_107_clock),
    .reset(FP_multiplier_10ccs_107_reset),
    .io_in_a(FP_multiplier_10ccs_107_io_in_a),
    .io_in_b(FP_multiplier_10ccs_107_io_in_b),
    .io_out_s(FP_multiplier_10ccs_107_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_108 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_108_clock),
    .reset(FP_multiplier_10ccs_108_reset),
    .io_in_a(FP_multiplier_10ccs_108_io_in_a),
    .io_in_b(FP_multiplier_10ccs_108_io_in_b),
    .io_out_s(FP_multiplier_10ccs_108_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_109 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_109_clock),
    .reset(FP_multiplier_10ccs_109_reset),
    .io_in_a(FP_multiplier_10ccs_109_io_in_a),
    .io_in_b(FP_multiplier_10ccs_109_io_in_b),
    .io_out_s(FP_multiplier_10ccs_109_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_110 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_110_clock),
    .reset(FP_multiplier_10ccs_110_reset),
    .io_in_a(FP_multiplier_10ccs_110_io_in_a),
    .io_in_b(FP_multiplier_10ccs_110_io_in_b),
    .io_out_s(FP_multiplier_10ccs_110_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_111 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_111_clock),
    .reset(FP_multiplier_10ccs_111_reset),
    .io_in_a(FP_multiplier_10ccs_111_io_in_a),
    .io_in_b(FP_multiplier_10ccs_111_io_in_b),
    .io_out_s(FP_multiplier_10ccs_111_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_112 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_112_clock),
    .reset(FP_multiplier_10ccs_112_reset),
    .io_in_a(FP_multiplier_10ccs_112_io_in_a),
    .io_in_b(FP_multiplier_10ccs_112_io_in_b),
    .io_out_s(FP_multiplier_10ccs_112_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_113 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_113_clock),
    .reset(FP_multiplier_10ccs_113_reset),
    .io_in_a(FP_multiplier_10ccs_113_io_in_a),
    .io_in_b(FP_multiplier_10ccs_113_io_in_b),
    .io_out_s(FP_multiplier_10ccs_113_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_114 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_114_clock),
    .reset(FP_multiplier_10ccs_114_reset),
    .io_in_a(FP_multiplier_10ccs_114_io_in_a),
    .io_in_b(FP_multiplier_10ccs_114_io_in_b),
    .io_out_s(FP_multiplier_10ccs_114_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_115 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_115_clock),
    .reset(FP_multiplier_10ccs_115_reset),
    .io_in_a(FP_multiplier_10ccs_115_io_in_a),
    .io_in_b(FP_multiplier_10ccs_115_io_in_b),
    .io_out_s(FP_multiplier_10ccs_115_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_116 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_116_clock),
    .reset(FP_multiplier_10ccs_116_reset),
    .io_in_a(FP_multiplier_10ccs_116_io_in_a),
    .io_in_b(FP_multiplier_10ccs_116_io_in_b),
    .io_out_s(FP_multiplier_10ccs_116_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_117 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_117_clock),
    .reset(FP_multiplier_10ccs_117_reset),
    .io_in_a(FP_multiplier_10ccs_117_io_in_a),
    .io_in_b(FP_multiplier_10ccs_117_io_in_b),
    .io_out_s(FP_multiplier_10ccs_117_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_118 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_118_clock),
    .reset(FP_multiplier_10ccs_118_reset),
    .io_in_a(FP_multiplier_10ccs_118_io_in_a),
    .io_in_b(FP_multiplier_10ccs_118_io_in_b),
    .io_out_s(FP_multiplier_10ccs_118_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_119 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_119_clock),
    .reset(FP_multiplier_10ccs_119_reset),
    .io_in_a(FP_multiplier_10ccs_119_io_in_a),
    .io_in_b(FP_multiplier_10ccs_119_io_in_b),
    .io_out_s(FP_multiplier_10ccs_119_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_120 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_120_clock),
    .reset(FP_multiplier_10ccs_120_reset),
    .io_in_a(FP_multiplier_10ccs_120_io_in_a),
    .io_in_b(FP_multiplier_10ccs_120_io_in_b),
    .io_out_s(FP_multiplier_10ccs_120_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_121 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_121_clock),
    .reset(FP_multiplier_10ccs_121_reset),
    .io_in_a(FP_multiplier_10ccs_121_io_in_a),
    .io_in_b(FP_multiplier_10ccs_121_io_in_b),
    .io_out_s(FP_multiplier_10ccs_121_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_122 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_122_clock),
    .reset(FP_multiplier_10ccs_122_reset),
    .io_in_a(FP_multiplier_10ccs_122_io_in_a),
    .io_in_b(FP_multiplier_10ccs_122_io_in_b),
    .io_out_s(FP_multiplier_10ccs_122_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_123 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_123_clock),
    .reset(FP_multiplier_10ccs_123_reset),
    .io_in_a(FP_multiplier_10ccs_123_io_in_a),
    .io_in_b(FP_multiplier_10ccs_123_io_in_b),
    .io_out_s(FP_multiplier_10ccs_123_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_124 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_124_clock),
    .reset(FP_multiplier_10ccs_124_reset),
    .io_in_a(FP_multiplier_10ccs_124_io_in_a),
    .io_in_b(FP_multiplier_10ccs_124_io_in_b),
    .io_out_s(FP_multiplier_10ccs_124_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_125 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_125_clock),
    .reset(FP_multiplier_10ccs_125_reset),
    .io_in_a(FP_multiplier_10ccs_125_io_in_a),
    .io_in_b(FP_multiplier_10ccs_125_io_in_b),
    .io_out_s(FP_multiplier_10ccs_125_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_126 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_126_clock),
    .reset(FP_multiplier_10ccs_126_reset),
    .io_in_a(FP_multiplier_10ccs_126_io_in_a),
    .io_in_b(FP_multiplier_10ccs_126_io_in_b),
    .io_out_s(FP_multiplier_10ccs_126_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_127 ( // @[FloatingPointDesigns.scala 2409:44]
    .clock(FP_multiplier_10ccs_127_clock),
    .reset(FP_multiplier_10ccs_127_reset),
    .io_in_a(FP_multiplier_10ccs_127_io_in_a),
    .io_in_b(FP_multiplier_10ccs_127_io_in_b),
    .io_out_s(FP_multiplier_10ccs_127_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_clock),
    .reset(FP_adder_13ccs_reset),
    .io_in_a(FP_adder_13ccs_io_in_a),
    .io_in_b(FP_adder_13ccs_io_in_b),
    .io_out_s(FP_adder_13ccs_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_1 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_1_clock),
    .reset(FP_adder_13ccs_1_reset),
    .io_in_a(FP_adder_13ccs_1_io_in_a),
    .io_in_b(FP_adder_13ccs_1_io_in_b),
    .io_out_s(FP_adder_13ccs_1_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_2 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_2_clock),
    .reset(FP_adder_13ccs_2_reset),
    .io_in_a(FP_adder_13ccs_2_io_in_a),
    .io_in_b(FP_adder_13ccs_2_io_in_b),
    .io_out_s(FP_adder_13ccs_2_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_3 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_3_clock),
    .reset(FP_adder_13ccs_3_reset),
    .io_in_a(FP_adder_13ccs_3_io_in_a),
    .io_in_b(FP_adder_13ccs_3_io_in_b),
    .io_out_s(FP_adder_13ccs_3_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_4 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_4_clock),
    .reset(FP_adder_13ccs_4_reset),
    .io_in_a(FP_adder_13ccs_4_io_in_a),
    .io_in_b(FP_adder_13ccs_4_io_in_b),
    .io_out_s(FP_adder_13ccs_4_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_5 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_5_clock),
    .reset(FP_adder_13ccs_5_reset),
    .io_in_a(FP_adder_13ccs_5_io_in_a),
    .io_in_b(FP_adder_13ccs_5_io_in_b),
    .io_out_s(FP_adder_13ccs_5_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_6 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_6_clock),
    .reset(FP_adder_13ccs_6_reset),
    .io_in_a(FP_adder_13ccs_6_io_in_a),
    .io_in_b(FP_adder_13ccs_6_io_in_b),
    .io_out_s(FP_adder_13ccs_6_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_7 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_7_clock),
    .reset(FP_adder_13ccs_7_reset),
    .io_in_a(FP_adder_13ccs_7_io_in_a),
    .io_in_b(FP_adder_13ccs_7_io_in_b),
    .io_out_s(FP_adder_13ccs_7_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_8 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_8_clock),
    .reset(FP_adder_13ccs_8_reset),
    .io_in_a(FP_adder_13ccs_8_io_in_a),
    .io_in_b(FP_adder_13ccs_8_io_in_b),
    .io_out_s(FP_adder_13ccs_8_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_9 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_9_clock),
    .reset(FP_adder_13ccs_9_reset),
    .io_in_a(FP_adder_13ccs_9_io_in_a),
    .io_in_b(FP_adder_13ccs_9_io_in_b),
    .io_out_s(FP_adder_13ccs_9_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_10 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_10_clock),
    .reset(FP_adder_13ccs_10_reset),
    .io_in_a(FP_adder_13ccs_10_io_in_a),
    .io_in_b(FP_adder_13ccs_10_io_in_b),
    .io_out_s(FP_adder_13ccs_10_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_11 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_11_clock),
    .reset(FP_adder_13ccs_11_reset),
    .io_in_a(FP_adder_13ccs_11_io_in_a),
    .io_in_b(FP_adder_13ccs_11_io_in_b),
    .io_out_s(FP_adder_13ccs_11_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_12 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_12_clock),
    .reset(FP_adder_13ccs_12_reset),
    .io_in_a(FP_adder_13ccs_12_io_in_a),
    .io_in_b(FP_adder_13ccs_12_io_in_b),
    .io_out_s(FP_adder_13ccs_12_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_13 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_13_clock),
    .reset(FP_adder_13ccs_13_reset),
    .io_in_a(FP_adder_13ccs_13_io_in_a),
    .io_in_b(FP_adder_13ccs_13_io_in_b),
    .io_out_s(FP_adder_13ccs_13_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_14 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_14_clock),
    .reset(FP_adder_13ccs_14_reset),
    .io_in_a(FP_adder_13ccs_14_io_in_a),
    .io_in_b(FP_adder_13ccs_14_io_in_b),
    .io_out_s(FP_adder_13ccs_14_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_15 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_15_clock),
    .reset(FP_adder_13ccs_15_reset),
    .io_in_a(FP_adder_13ccs_15_io_in_a),
    .io_in_b(FP_adder_13ccs_15_io_in_b),
    .io_out_s(FP_adder_13ccs_15_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_16 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_16_clock),
    .reset(FP_adder_13ccs_16_reset),
    .io_in_a(FP_adder_13ccs_16_io_in_a),
    .io_in_b(FP_adder_13ccs_16_io_in_b),
    .io_out_s(FP_adder_13ccs_16_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_17 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_17_clock),
    .reset(FP_adder_13ccs_17_reset),
    .io_in_a(FP_adder_13ccs_17_io_in_a),
    .io_in_b(FP_adder_13ccs_17_io_in_b),
    .io_out_s(FP_adder_13ccs_17_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_18 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_18_clock),
    .reset(FP_adder_13ccs_18_reset),
    .io_in_a(FP_adder_13ccs_18_io_in_a),
    .io_in_b(FP_adder_13ccs_18_io_in_b),
    .io_out_s(FP_adder_13ccs_18_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_19 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_19_clock),
    .reset(FP_adder_13ccs_19_reset),
    .io_in_a(FP_adder_13ccs_19_io_in_a),
    .io_in_b(FP_adder_13ccs_19_io_in_b),
    .io_out_s(FP_adder_13ccs_19_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_20 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_20_clock),
    .reset(FP_adder_13ccs_20_reset),
    .io_in_a(FP_adder_13ccs_20_io_in_a),
    .io_in_b(FP_adder_13ccs_20_io_in_b),
    .io_out_s(FP_adder_13ccs_20_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_21 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_21_clock),
    .reset(FP_adder_13ccs_21_reset),
    .io_in_a(FP_adder_13ccs_21_io_in_a),
    .io_in_b(FP_adder_13ccs_21_io_in_b),
    .io_out_s(FP_adder_13ccs_21_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_22 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_22_clock),
    .reset(FP_adder_13ccs_22_reset),
    .io_in_a(FP_adder_13ccs_22_io_in_a),
    .io_in_b(FP_adder_13ccs_22_io_in_b),
    .io_out_s(FP_adder_13ccs_22_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_23 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_23_clock),
    .reset(FP_adder_13ccs_23_reset),
    .io_in_a(FP_adder_13ccs_23_io_in_a),
    .io_in_b(FP_adder_13ccs_23_io_in_b),
    .io_out_s(FP_adder_13ccs_23_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_24 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_24_clock),
    .reset(FP_adder_13ccs_24_reset),
    .io_in_a(FP_adder_13ccs_24_io_in_a),
    .io_in_b(FP_adder_13ccs_24_io_in_b),
    .io_out_s(FP_adder_13ccs_24_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_25 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_25_clock),
    .reset(FP_adder_13ccs_25_reset),
    .io_in_a(FP_adder_13ccs_25_io_in_a),
    .io_in_b(FP_adder_13ccs_25_io_in_b),
    .io_out_s(FP_adder_13ccs_25_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_26 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_26_clock),
    .reset(FP_adder_13ccs_26_reset),
    .io_in_a(FP_adder_13ccs_26_io_in_a),
    .io_in_b(FP_adder_13ccs_26_io_in_b),
    .io_out_s(FP_adder_13ccs_26_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_27 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_27_clock),
    .reset(FP_adder_13ccs_27_reset),
    .io_in_a(FP_adder_13ccs_27_io_in_a),
    .io_in_b(FP_adder_13ccs_27_io_in_b),
    .io_out_s(FP_adder_13ccs_27_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_28 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_28_clock),
    .reset(FP_adder_13ccs_28_reset),
    .io_in_a(FP_adder_13ccs_28_io_in_a),
    .io_in_b(FP_adder_13ccs_28_io_in_b),
    .io_out_s(FP_adder_13ccs_28_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_29 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_29_clock),
    .reset(FP_adder_13ccs_29_reset),
    .io_in_a(FP_adder_13ccs_29_io_in_a),
    .io_in_b(FP_adder_13ccs_29_io_in_b),
    .io_out_s(FP_adder_13ccs_29_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_30 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_30_clock),
    .reset(FP_adder_13ccs_30_reset),
    .io_in_a(FP_adder_13ccs_30_io_in_a),
    .io_in_b(FP_adder_13ccs_30_io_in_b),
    .io_out_s(FP_adder_13ccs_30_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_31 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_31_clock),
    .reset(FP_adder_13ccs_31_reset),
    .io_in_a(FP_adder_13ccs_31_io_in_a),
    .io_in_b(FP_adder_13ccs_31_io_in_b),
    .io_out_s(FP_adder_13ccs_31_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_32 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_32_clock),
    .reset(FP_adder_13ccs_32_reset),
    .io_in_a(FP_adder_13ccs_32_io_in_a),
    .io_in_b(FP_adder_13ccs_32_io_in_b),
    .io_out_s(FP_adder_13ccs_32_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_33 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_33_clock),
    .reset(FP_adder_13ccs_33_reset),
    .io_in_a(FP_adder_13ccs_33_io_in_a),
    .io_in_b(FP_adder_13ccs_33_io_in_b),
    .io_out_s(FP_adder_13ccs_33_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_34 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_34_clock),
    .reset(FP_adder_13ccs_34_reset),
    .io_in_a(FP_adder_13ccs_34_io_in_a),
    .io_in_b(FP_adder_13ccs_34_io_in_b),
    .io_out_s(FP_adder_13ccs_34_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_35 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_35_clock),
    .reset(FP_adder_13ccs_35_reset),
    .io_in_a(FP_adder_13ccs_35_io_in_a),
    .io_in_b(FP_adder_13ccs_35_io_in_b),
    .io_out_s(FP_adder_13ccs_35_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_36 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_36_clock),
    .reset(FP_adder_13ccs_36_reset),
    .io_in_a(FP_adder_13ccs_36_io_in_a),
    .io_in_b(FP_adder_13ccs_36_io_in_b),
    .io_out_s(FP_adder_13ccs_36_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_37 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_37_clock),
    .reset(FP_adder_13ccs_37_reset),
    .io_in_a(FP_adder_13ccs_37_io_in_a),
    .io_in_b(FP_adder_13ccs_37_io_in_b),
    .io_out_s(FP_adder_13ccs_37_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_38 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_38_clock),
    .reset(FP_adder_13ccs_38_reset),
    .io_in_a(FP_adder_13ccs_38_io_in_a),
    .io_in_b(FP_adder_13ccs_38_io_in_b),
    .io_out_s(FP_adder_13ccs_38_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_39 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_39_clock),
    .reset(FP_adder_13ccs_39_reset),
    .io_in_a(FP_adder_13ccs_39_io_in_a),
    .io_in_b(FP_adder_13ccs_39_io_in_b),
    .io_out_s(FP_adder_13ccs_39_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_40 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_40_clock),
    .reset(FP_adder_13ccs_40_reset),
    .io_in_a(FP_adder_13ccs_40_io_in_a),
    .io_in_b(FP_adder_13ccs_40_io_in_b),
    .io_out_s(FP_adder_13ccs_40_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_41 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_41_clock),
    .reset(FP_adder_13ccs_41_reset),
    .io_in_a(FP_adder_13ccs_41_io_in_a),
    .io_in_b(FP_adder_13ccs_41_io_in_b),
    .io_out_s(FP_adder_13ccs_41_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_42 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_42_clock),
    .reset(FP_adder_13ccs_42_reset),
    .io_in_a(FP_adder_13ccs_42_io_in_a),
    .io_in_b(FP_adder_13ccs_42_io_in_b),
    .io_out_s(FP_adder_13ccs_42_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_43 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_43_clock),
    .reset(FP_adder_13ccs_43_reset),
    .io_in_a(FP_adder_13ccs_43_io_in_a),
    .io_in_b(FP_adder_13ccs_43_io_in_b),
    .io_out_s(FP_adder_13ccs_43_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_44 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_44_clock),
    .reset(FP_adder_13ccs_44_reset),
    .io_in_a(FP_adder_13ccs_44_io_in_a),
    .io_in_b(FP_adder_13ccs_44_io_in_b),
    .io_out_s(FP_adder_13ccs_44_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_45 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_45_clock),
    .reset(FP_adder_13ccs_45_reset),
    .io_in_a(FP_adder_13ccs_45_io_in_a),
    .io_in_b(FP_adder_13ccs_45_io_in_b),
    .io_out_s(FP_adder_13ccs_45_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_46 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_46_clock),
    .reset(FP_adder_13ccs_46_reset),
    .io_in_a(FP_adder_13ccs_46_io_in_a),
    .io_in_b(FP_adder_13ccs_46_io_in_b),
    .io_out_s(FP_adder_13ccs_46_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_47 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_47_clock),
    .reset(FP_adder_13ccs_47_reset),
    .io_in_a(FP_adder_13ccs_47_io_in_a),
    .io_in_b(FP_adder_13ccs_47_io_in_b),
    .io_out_s(FP_adder_13ccs_47_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_48 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_48_clock),
    .reset(FP_adder_13ccs_48_reset),
    .io_in_a(FP_adder_13ccs_48_io_in_a),
    .io_in_b(FP_adder_13ccs_48_io_in_b),
    .io_out_s(FP_adder_13ccs_48_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_49 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_49_clock),
    .reset(FP_adder_13ccs_49_reset),
    .io_in_a(FP_adder_13ccs_49_io_in_a),
    .io_in_b(FP_adder_13ccs_49_io_in_b),
    .io_out_s(FP_adder_13ccs_49_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_50 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_50_clock),
    .reset(FP_adder_13ccs_50_reset),
    .io_in_a(FP_adder_13ccs_50_io_in_a),
    .io_in_b(FP_adder_13ccs_50_io_in_b),
    .io_out_s(FP_adder_13ccs_50_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_51 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_51_clock),
    .reset(FP_adder_13ccs_51_reset),
    .io_in_a(FP_adder_13ccs_51_io_in_a),
    .io_in_b(FP_adder_13ccs_51_io_in_b),
    .io_out_s(FP_adder_13ccs_51_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_52 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_52_clock),
    .reset(FP_adder_13ccs_52_reset),
    .io_in_a(FP_adder_13ccs_52_io_in_a),
    .io_in_b(FP_adder_13ccs_52_io_in_b),
    .io_out_s(FP_adder_13ccs_52_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_53 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_53_clock),
    .reset(FP_adder_13ccs_53_reset),
    .io_in_a(FP_adder_13ccs_53_io_in_a),
    .io_in_b(FP_adder_13ccs_53_io_in_b),
    .io_out_s(FP_adder_13ccs_53_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_54 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_54_clock),
    .reset(FP_adder_13ccs_54_reset),
    .io_in_a(FP_adder_13ccs_54_io_in_a),
    .io_in_b(FP_adder_13ccs_54_io_in_b),
    .io_out_s(FP_adder_13ccs_54_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_55 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_55_clock),
    .reset(FP_adder_13ccs_55_reset),
    .io_in_a(FP_adder_13ccs_55_io_in_a),
    .io_in_b(FP_adder_13ccs_55_io_in_b),
    .io_out_s(FP_adder_13ccs_55_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_56 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_56_clock),
    .reset(FP_adder_13ccs_56_reset),
    .io_in_a(FP_adder_13ccs_56_io_in_a),
    .io_in_b(FP_adder_13ccs_56_io_in_b),
    .io_out_s(FP_adder_13ccs_56_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_57 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_57_clock),
    .reset(FP_adder_13ccs_57_reset),
    .io_in_a(FP_adder_13ccs_57_io_in_a),
    .io_in_b(FP_adder_13ccs_57_io_in_b),
    .io_out_s(FP_adder_13ccs_57_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_58 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_58_clock),
    .reset(FP_adder_13ccs_58_reset),
    .io_in_a(FP_adder_13ccs_58_io_in_a),
    .io_in_b(FP_adder_13ccs_58_io_in_b),
    .io_out_s(FP_adder_13ccs_58_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_59 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_59_clock),
    .reset(FP_adder_13ccs_59_reset),
    .io_in_a(FP_adder_13ccs_59_io_in_a),
    .io_in_b(FP_adder_13ccs_59_io_in_b),
    .io_out_s(FP_adder_13ccs_59_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_60 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_60_clock),
    .reset(FP_adder_13ccs_60_reset),
    .io_in_a(FP_adder_13ccs_60_io_in_a),
    .io_in_b(FP_adder_13ccs_60_io_in_b),
    .io_out_s(FP_adder_13ccs_60_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_61 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_61_clock),
    .reset(FP_adder_13ccs_61_reset),
    .io_in_a(FP_adder_13ccs_61_io_in_a),
    .io_in_b(FP_adder_13ccs_61_io_in_b),
    .io_out_s(FP_adder_13ccs_61_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_62 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_62_clock),
    .reset(FP_adder_13ccs_62_reset),
    .io_in_a(FP_adder_13ccs_62_io_in_a),
    .io_in_b(FP_adder_13ccs_62_io_in_b),
    .io_out_s(FP_adder_13ccs_62_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_63 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_63_clock),
    .reset(FP_adder_13ccs_63_reset),
    .io_in_a(FP_adder_13ccs_63_io_in_a),
    .io_in_b(FP_adder_13ccs_63_io_in_b),
    .io_out_s(FP_adder_13ccs_63_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_64 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_64_clock),
    .reset(FP_adder_13ccs_64_reset),
    .io_in_a(FP_adder_13ccs_64_io_in_a),
    .io_in_b(FP_adder_13ccs_64_io_in_b),
    .io_out_s(FP_adder_13ccs_64_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_65 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_65_clock),
    .reset(FP_adder_13ccs_65_reset),
    .io_in_a(FP_adder_13ccs_65_io_in_a),
    .io_in_b(FP_adder_13ccs_65_io_in_b),
    .io_out_s(FP_adder_13ccs_65_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_66 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_66_clock),
    .reset(FP_adder_13ccs_66_reset),
    .io_in_a(FP_adder_13ccs_66_io_in_a),
    .io_in_b(FP_adder_13ccs_66_io_in_b),
    .io_out_s(FP_adder_13ccs_66_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_67 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_67_clock),
    .reset(FP_adder_13ccs_67_reset),
    .io_in_a(FP_adder_13ccs_67_io_in_a),
    .io_in_b(FP_adder_13ccs_67_io_in_b),
    .io_out_s(FP_adder_13ccs_67_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_68 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_68_clock),
    .reset(FP_adder_13ccs_68_reset),
    .io_in_a(FP_adder_13ccs_68_io_in_a),
    .io_in_b(FP_adder_13ccs_68_io_in_b),
    .io_out_s(FP_adder_13ccs_68_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_69 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_69_clock),
    .reset(FP_adder_13ccs_69_reset),
    .io_in_a(FP_adder_13ccs_69_io_in_a),
    .io_in_b(FP_adder_13ccs_69_io_in_b),
    .io_out_s(FP_adder_13ccs_69_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_70 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_70_clock),
    .reset(FP_adder_13ccs_70_reset),
    .io_in_a(FP_adder_13ccs_70_io_in_a),
    .io_in_b(FP_adder_13ccs_70_io_in_b),
    .io_out_s(FP_adder_13ccs_70_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_71 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_71_clock),
    .reset(FP_adder_13ccs_71_reset),
    .io_in_a(FP_adder_13ccs_71_io_in_a),
    .io_in_b(FP_adder_13ccs_71_io_in_b),
    .io_out_s(FP_adder_13ccs_71_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_72 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_72_clock),
    .reset(FP_adder_13ccs_72_reset),
    .io_in_a(FP_adder_13ccs_72_io_in_a),
    .io_in_b(FP_adder_13ccs_72_io_in_b),
    .io_out_s(FP_adder_13ccs_72_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_73 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_73_clock),
    .reset(FP_adder_13ccs_73_reset),
    .io_in_a(FP_adder_13ccs_73_io_in_a),
    .io_in_b(FP_adder_13ccs_73_io_in_b),
    .io_out_s(FP_adder_13ccs_73_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_74 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_74_clock),
    .reset(FP_adder_13ccs_74_reset),
    .io_in_a(FP_adder_13ccs_74_io_in_a),
    .io_in_b(FP_adder_13ccs_74_io_in_b),
    .io_out_s(FP_adder_13ccs_74_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_75 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_75_clock),
    .reset(FP_adder_13ccs_75_reset),
    .io_in_a(FP_adder_13ccs_75_io_in_a),
    .io_in_b(FP_adder_13ccs_75_io_in_b),
    .io_out_s(FP_adder_13ccs_75_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_76 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_76_clock),
    .reset(FP_adder_13ccs_76_reset),
    .io_in_a(FP_adder_13ccs_76_io_in_a),
    .io_in_b(FP_adder_13ccs_76_io_in_b),
    .io_out_s(FP_adder_13ccs_76_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_77 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_77_clock),
    .reset(FP_adder_13ccs_77_reset),
    .io_in_a(FP_adder_13ccs_77_io_in_a),
    .io_in_b(FP_adder_13ccs_77_io_in_b),
    .io_out_s(FP_adder_13ccs_77_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_78 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_78_clock),
    .reset(FP_adder_13ccs_78_reset),
    .io_in_a(FP_adder_13ccs_78_io_in_a),
    .io_in_b(FP_adder_13ccs_78_io_in_b),
    .io_out_s(FP_adder_13ccs_78_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_79 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_79_clock),
    .reset(FP_adder_13ccs_79_reset),
    .io_in_a(FP_adder_13ccs_79_io_in_a),
    .io_in_b(FP_adder_13ccs_79_io_in_b),
    .io_out_s(FP_adder_13ccs_79_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_80 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_80_clock),
    .reset(FP_adder_13ccs_80_reset),
    .io_in_a(FP_adder_13ccs_80_io_in_a),
    .io_in_b(FP_adder_13ccs_80_io_in_b),
    .io_out_s(FP_adder_13ccs_80_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_81 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_81_clock),
    .reset(FP_adder_13ccs_81_reset),
    .io_in_a(FP_adder_13ccs_81_io_in_a),
    .io_in_b(FP_adder_13ccs_81_io_in_b),
    .io_out_s(FP_adder_13ccs_81_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_82 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_82_clock),
    .reset(FP_adder_13ccs_82_reset),
    .io_in_a(FP_adder_13ccs_82_io_in_a),
    .io_in_b(FP_adder_13ccs_82_io_in_b),
    .io_out_s(FP_adder_13ccs_82_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_83 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_83_clock),
    .reset(FP_adder_13ccs_83_reset),
    .io_in_a(FP_adder_13ccs_83_io_in_a),
    .io_in_b(FP_adder_13ccs_83_io_in_b),
    .io_out_s(FP_adder_13ccs_83_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_84 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_84_clock),
    .reset(FP_adder_13ccs_84_reset),
    .io_in_a(FP_adder_13ccs_84_io_in_a),
    .io_in_b(FP_adder_13ccs_84_io_in_b),
    .io_out_s(FP_adder_13ccs_84_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_85 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_85_clock),
    .reset(FP_adder_13ccs_85_reset),
    .io_in_a(FP_adder_13ccs_85_io_in_a),
    .io_in_b(FP_adder_13ccs_85_io_in_b),
    .io_out_s(FP_adder_13ccs_85_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_86 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_86_clock),
    .reset(FP_adder_13ccs_86_reset),
    .io_in_a(FP_adder_13ccs_86_io_in_a),
    .io_in_b(FP_adder_13ccs_86_io_in_b),
    .io_out_s(FP_adder_13ccs_86_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_87 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_87_clock),
    .reset(FP_adder_13ccs_87_reset),
    .io_in_a(FP_adder_13ccs_87_io_in_a),
    .io_in_b(FP_adder_13ccs_87_io_in_b),
    .io_out_s(FP_adder_13ccs_87_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_88 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_88_clock),
    .reset(FP_adder_13ccs_88_reset),
    .io_in_a(FP_adder_13ccs_88_io_in_a),
    .io_in_b(FP_adder_13ccs_88_io_in_b),
    .io_out_s(FP_adder_13ccs_88_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_89 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_89_clock),
    .reset(FP_adder_13ccs_89_reset),
    .io_in_a(FP_adder_13ccs_89_io_in_a),
    .io_in_b(FP_adder_13ccs_89_io_in_b),
    .io_out_s(FP_adder_13ccs_89_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_90 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_90_clock),
    .reset(FP_adder_13ccs_90_reset),
    .io_in_a(FP_adder_13ccs_90_io_in_a),
    .io_in_b(FP_adder_13ccs_90_io_in_b),
    .io_out_s(FP_adder_13ccs_90_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_91 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_91_clock),
    .reset(FP_adder_13ccs_91_reset),
    .io_in_a(FP_adder_13ccs_91_io_in_a),
    .io_in_b(FP_adder_13ccs_91_io_in_b),
    .io_out_s(FP_adder_13ccs_91_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_92 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_92_clock),
    .reset(FP_adder_13ccs_92_reset),
    .io_in_a(FP_adder_13ccs_92_io_in_a),
    .io_in_b(FP_adder_13ccs_92_io_in_b),
    .io_out_s(FP_adder_13ccs_92_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_93 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_93_clock),
    .reset(FP_adder_13ccs_93_reset),
    .io_in_a(FP_adder_13ccs_93_io_in_a),
    .io_in_b(FP_adder_13ccs_93_io_in_b),
    .io_out_s(FP_adder_13ccs_93_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_94 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_94_clock),
    .reset(FP_adder_13ccs_94_reset),
    .io_in_a(FP_adder_13ccs_94_io_in_a),
    .io_in_b(FP_adder_13ccs_94_io_in_b),
    .io_out_s(FP_adder_13ccs_94_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_95 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_95_clock),
    .reset(FP_adder_13ccs_95_reset),
    .io_in_a(FP_adder_13ccs_95_io_in_a),
    .io_in_b(FP_adder_13ccs_95_io_in_b),
    .io_out_s(FP_adder_13ccs_95_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_96 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_96_clock),
    .reset(FP_adder_13ccs_96_reset),
    .io_in_a(FP_adder_13ccs_96_io_in_a),
    .io_in_b(FP_adder_13ccs_96_io_in_b),
    .io_out_s(FP_adder_13ccs_96_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_97 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_97_clock),
    .reset(FP_adder_13ccs_97_reset),
    .io_in_a(FP_adder_13ccs_97_io_in_a),
    .io_in_b(FP_adder_13ccs_97_io_in_b),
    .io_out_s(FP_adder_13ccs_97_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_98 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_98_clock),
    .reset(FP_adder_13ccs_98_reset),
    .io_in_a(FP_adder_13ccs_98_io_in_a),
    .io_in_b(FP_adder_13ccs_98_io_in_b),
    .io_out_s(FP_adder_13ccs_98_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_99 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_99_clock),
    .reset(FP_adder_13ccs_99_reset),
    .io_in_a(FP_adder_13ccs_99_io_in_a),
    .io_in_b(FP_adder_13ccs_99_io_in_b),
    .io_out_s(FP_adder_13ccs_99_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_100 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_100_clock),
    .reset(FP_adder_13ccs_100_reset),
    .io_in_a(FP_adder_13ccs_100_io_in_a),
    .io_in_b(FP_adder_13ccs_100_io_in_b),
    .io_out_s(FP_adder_13ccs_100_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_101 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_101_clock),
    .reset(FP_adder_13ccs_101_reset),
    .io_in_a(FP_adder_13ccs_101_io_in_a),
    .io_in_b(FP_adder_13ccs_101_io_in_b),
    .io_out_s(FP_adder_13ccs_101_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_102 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_102_clock),
    .reset(FP_adder_13ccs_102_reset),
    .io_in_a(FP_adder_13ccs_102_io_in_a),
    .io_in_b(FP_adder_13ccs_102_io_in_b),
    .io_out_s(FP_adder_13ccs_102_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_103 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_103_clock),
    .reset(FP_adder_13ccs_103_reset),
    .io_in_a(FP_adder_13ccs_103_io_in_a),
    .io_in_b(FP_adder_13ccs_103_io_in_b),
    .io_out_s(FP_adder_13ccs_103_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_104 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_104_clock),
    .reset(FP_adder_13ccs_104_reset),
    .io_in_a(FP_adder_13ccs_104_io_in_a),
    .io_in_b(FP_adder_13ccs_104_io_in_b),
    .io_out_s(FP_adder_13ccs_104_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_105 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_105_clock),
    .reset(FP_adder_13ccs_105_reset),
    .io_in_a(FP_adder_13ccs_105_io_in_a),
    .io_in_b(FP_adder_13ccs_105_io_in_b),
    .io_out_s(FP_adder_13ccs_105_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_106 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_106_clock),
    .reset(FP_adder_13ccs_106_reset),
    .io_in_a(FP_adder_13ccs_106_io_in_a),
    .io_in_b(FP_adder_13ccs_106_io_in_b),
    .io_out_s(FP_adder_13ccs_106_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_107 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_107_clock),
    .reset(FP_adder_13ccs_107_reset),
    .io_in_a(FP_adder_13ccs_107_io_in_a),
    .io_in_b(FP_adder_13ccs_107_io_in_b),
    .io_out_s(FP_adder_13ccs_107_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_108 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_108_clock),
    .reset(FP_adder_13ccs_108_reset),
    .io_in_a(FP_adder_13ccs_108_io_in_a),
    .io_in_b(FP_adder_13ccs_108_io_in_b),
    .io_out_s(FP_adder_13ccs_108_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_109 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_109_clock),
    .reset(FP_adder_13ccs_109_reset),
    .io_in_a(FP_adder_13ccs_109_io_in_a),
    .io_in_b(FP_adder_13ccs_109_io_in_b),
    .io_out_s(FP_adder_13ccs_109_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_110 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_110_clock),
    .reset(FP_adder_13ccs_110_reset),
    .io_in_a(FP_adder_13ccs_110_io_in_a),
    .io_in_b(FP_adder_13ccs_110_io_in_b),
    .io_out_s(FP_adder_13ccs_110_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_111 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_111_clock),
    .reset(FP_adder_13ccs_111_reset),
    .io_in_a(FP_adder_13ccs_111_io_in_a),
    .io_in_b(FP_adder_13ccs_111_io_in_b),
    .io_out_s(FP_adder_13ccs_111_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_112 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_112_clock),
    .reset(FP_adder_13ccs_112_reset),
    .io_in_a(FP_adder_13ccs_112_io_in_a),
    .io_in_b(FP_adder_13ccs_112_io_in_b),
    .io_out_s(FP_adder_13ccs_112_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_113 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_113_clock),
    .reset(FP_adder_13ccs_113_reset),
    .io_in_a(FP_adder_13ccs_113_io_in_a),
    .io_in_b(FP_adder_13ccs_113_io_in_b),
    .io_out_s(FP_adder_13ccs_113_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_114 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_114_clock),
    .reset(FP_adder_13ccs_114_reset),
    .io_in_a(FP_adder_13ccs_114_io_in_a),
    .io_in_b(FP_adder_13ccs_114_io_in_b),
    .io_out_s(FP_adder_13ccs_114_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_115 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_115_clock),
    .reset(FP_adder_13ccs_115_reset),
    .io_in_a(FP_adder_13ccs_115_io_in_a),
    .io_in_b(FP_adder_13ccs_115_io_in_b),
    .io_out_s(FP_adder_13ccs_115_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_116 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_116_clock),
    .reset(FP_adder_13ccs_116_reset),
    .io_in_a(FP_adder_13ccs_116_io_in_a),
    .io_in_b(FP_adder_13ccs_116_io_in_b),
    .io_out_s(FP_adder_13ccs_116_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_117 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_117_clock),
    .reset(FP_adder_13ccs_117_reset),
    .io_in_a(FP_adder_13ccs_117_io_in_a),
    .io_in_b(FP_adder_13ccs_117_io_in_b),
    .io_out_s(FP_adder_13ccs_117_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_118 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_118_clock),
    .reset(FP_adder_13ccs_118_reset),
    .io_in_a(FP_adder_13ccs_118_io_in_a),
    .io_in_b(FP_adder_13ccs_118_io_in_b),
    .io_out_s(FP_adder_13ccs_118_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_119 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_119_clock),
    .reset(FP_adder_13ccs_119_reset),
    .io_in_a(FP_adder_13ccs_119_io_in_a),
    .io_in_b(FP_adder_13ccs_119_io_in_b),
    .io_out_s(FP_adder_13ccs_119_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_120 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_120_clock),
    .reset(FP_adder_13ccs_120_reset),
    .io_in_a(FP_adder_13ccs_120_io_in_a),
    .io_in_b(FP_adder_13ccs_120_io_in_b),
    .io_out_s(FP_adder_13ccs_120_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_121 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_121_clock),
    .reset(FP_adder_13ccs_121_reset),
    .io_in_a(FP_adder_13ccs_121_io_in_a),
    .io_in_b(FP_adder_13ccs_121_io_in_b),
    .io_out_s(FP_adder_13ccs_121_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_122 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_122_clock),
    .reset(FP_adder_13ccs_122_reset),
    .io_in_a(FP_adder_13ccs_122_io_in_a),
    .io_in_b(FP_adder_13ccs_122_io_in_b),
    .io_out_s(FP_adder_13ccs_122_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_123 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_123_clock),
    .reset(FP_adder_13ccs_123_reset),
    .io_in_a(FP_adder_13ccs_123_io_in_a),
    .io_in_b(FP_adder_13ccs_123_io_in_b),
    .io_out_s(FP_adder_13ccs_123_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_124 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_124_clock),
    .reset(FP_adder_13ccs_124_reset),
    .io_in_a(FP_adder_13ccs_124_io_in_a),
    .io_in_b(FP_adder_13ccs_124_io_in_b),
    .io_out_s(FP_adder_13ccs_124_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_125 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_125_clock),
    .reset(FP_adder_13ccs_125_reset),
    .io_in_a(FP_adder_13ccs_125_io_in_a),
    .io_in_b(FP_adder_13ccs_125_io_in_b),
    .io_out_s(FP_adder_13ccs_125_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_126 ( // @[FloatingPointDesigns.scala 2417:17]
    .clock(FP_adder_13ccs_126_clock),
    .reset(FP_adder_13ccs_126_reset),
    .io_in_a(FP_adder_13ccs_126_io_in_a),
    .io_in_b(FP_adder_13ccs_126_io_in_b),
    .io_out_s(FP_adder_13ccs_126_io_out_s)
  );
  assign io_out_s = FP_adder_13ccs_126_io_out_s; // @[FloatingPointDesigns.scala 2466:16]
  assign FP_multiplier_10ccs_clock = clock;
  assign FP_multiplier_10ccs_reset = reset;
  assign FP_multiplier_10ccs_io_in_a = io_in_a_0; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_io_in_b = io_in_b_0; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_1_clock = clock;
  assign FP_multiplier_10ccs_1_reset = reset;
  assign FP_multiplier_10ccs_1_io_in_a = io_in_a_1; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_1_io_in_b = io_in_b_1; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_2_clock = clock;
  assign FP_multiplier_10ccs_2_reset = reset;
  assign FP_multiplier_10ccs_2_io_in_a = io_in_a_2; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_2_io_in_b = io_in_b_2; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_3_clock = clock;
  assign FP_multiplier_10ccs_3_reset = reset;
  assign FP_multiplier_10ccs_3_io_in_a = io_in_a_3; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_3_io_in_b = io_in_b_3; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_4_clock = clock;
  assign FP_multiplier_10ccs_4_reset = reset;
  assign FP_multiplier_10ccs_4_io_in_a = io_in_a_4; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_4_io_in_b = io_in_b_4; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_5_clock = clock;
  assign FP_multiplier_10ccs_5_reset = reset;
  assign FP_multiplier_10ccs_5_io_in_a = io_in_a_5; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_5_io_in_b = io_in_b_5; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_6_clock = clock;
  assign FP_multiplier_10ccs_6_reset = reset;
  assign FP_multiplier_10ccs_6_io_in_a = io_in_a_6; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_6_io_in_b = io_in_b_6; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_7_clock = clock;
  assign FP_multiplier_10ccs_7_reset = reset;
  assign FP_multiplier_10ccs_7_io_in_a = io_in_a_7; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_7_io_in_b = io_in_b_7; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_8_clock = clock;
  assign FP_multiplier_10ccs_8_reset = reset;
  assign FP_multiplier_10ccs_8_io_in_a = io_in_a_8; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_8_io_in_b = io_in_b_8; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_9_clock = clock;
  assign FP_multiplier_10ccs_9_reset = reset;
  assign FP_multiplier_10ccs_9_io_in_a = io_in_a_9; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_9_io_in_b = io_in_b_9; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_10_clock = clock;
  assign FP_multiplier_10ccs_10_reset = reset;
  assign FP_multiplier_10ccs_10_io_in_a = io_in_a_10; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_10_io_in_b = io_in_b_10; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_11_clock = clock;
  assign FP_multiplier_10ccs_11_reset = reset;
  assign FP_multiplier_10ccs_11_io_in_a = io_in_a_11; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_11_io_in_b = io_in_b_11; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_12_clock = clock;
  assign FP_multiplier_10ccs_12_reset = reset;
  assign FP_multiplier_10ccs_12_io_in_a = io_in_a_12; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_12_io_in_b = io_in_b_12; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_13_clock = clock;
  assign FP_multiplier_10ccs_13_reset = reset;
  assign FP_multiplier_10ccs_13_io_in_a = io_in_a_13; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_13_io_in_b = io_in_b_13; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_14_clock = clock;
  assign FP_multiplier_10ccs_14_reset = reset;
  assign FP_multiplier_10ccs_14_io_in_a = io_in_a_14; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_14_io_in_b = io_in_b_14; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_15_clock = clock;
  assign FP_multiplier_10ccs_15_reset = reset;
  assign FP_multiplier_10ccs_15_io_in_a = io_in_a_15; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_15_io_in_b = io_in_b_15; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_16_clock = clock;
  assign FP_multiplier_10ccs_16_reset = reset;
  assign FP_multiplier_10ccs_16_io_in_a = io_in_a_16; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_16_io_in_b = io_in_b_16; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_17_clock = clock;
  assign FP_multiplier_10ccs_17_reset = reset;
  assign FP_multiplier_10ccs_17_io_in_a = io_in_a_17; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_17_io_in_b = io_in_b_17; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_18_clock = clock;
  assign FP_multiplier_10ccs_18_reset = reset;
  assign FP_multiplier_10ccs_18_io_in_a = io_in_a_18; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_18_io_in_b = io_in_b_18; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_19_clock = clock;
  assign FP_multiplier_10ccs_19_reset = reset;
  assign FP_multiplier_10ccs_19_io_in_a = io_in_a_19; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_19_io_in_b = io_in_b_19; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_20_clock = clock;
  assign FP_multiplier_10ccs_20_reset = reset;
  assign FP_multiplier_10ccs_20_io_in_a = io_in_a_20; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_20_io_in_b = io_in_b_20; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_21_clock = clock;
  assign FP_multiplier_10ccs_21_reset = reset;
  assign FP_multiplier_10ccs_21_io_in_a = io_in_a_21; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_21_io_in_b = io_in_b_21; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_22_clock = clock;
  assign FP_multiplier_10ccs_22_reset = reset;
  assign FP_multiplier_10ccs_22_io_in_a = io_in_a_22; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_22_io_in_b = io_in_b_22; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_23_clock = clock;
  assign FP_multiplier_10ccs_23_reset = reset;
  assign FP_multiplier_10ccs_23_io_in_a = io_in_a_23; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_23_io_in_b = io_in_b_23; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_24_clock = clock;
  assign FP_multiplier_10ccs_24_reset = reset;
  assign FP_multiplier_10ccs_24_io_in_a = io_in_a_24; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_24_io_in_b = io_in_b_24; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_25_clock = clock;
  assign FP_multiplier_10ccs_25_reset = reset;
  assign FP_multiplier_10ccs_25_io_in_a = io_in_a_25; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_25_io_in_b = io_in_b_25; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_26_clock = clock;
  assign FP_multiplier_10ccs_26_reset = reset;
  assign FP_multiplier_10ccs_26_io_in_a = io_in_a_26; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_26_io_in_b = io_in_b_26; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_27_clock = clock;
  assign FP_multiplier_10ccs_27_reset = reset;
  assign FP_multiplier_10ccs_27_io_in_a = io_in_a_27; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_27_io_in_b = io_in_b_27; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_28_clock = clock;
  assign FP_multiplier_10ccs_28_reset = reset;
  assign FP_multiplier_10ccs_28_io_in_a = io_in_a_28; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_28_io_in_b = io_in_b_28; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_29_clock = clock;
  assign FP_multiplier_10ccs_29_reset = reset;
  assign FP_multiplier_10ccs_29_io_in_a = io_in_a_29; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_29_io_in_b = io_in_b_29; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_30_clock = clock;
  assign FP_multiplier_10ccs_30_reset = reset;
  assign FP_multiplier_10ccs_30_io_in_a = io_in_a_30; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_30_io_in_b = io_in_b_30; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_31_clock = clock;
  assign FP_multiplier_10ccs_31_reset = reset;
  assign FP_multiplier_10ccs_31_io_in_a = io_in_a_31; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_31_io_in_b = io_in_b_31; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_32_clock = clock;
  assign FP_multiplier_10ccs_32_reset = reset;
  assign FP_multiplier_10ccs_32_io_in_a = io_in_a_32; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_32_io_in_b = io_in_b_32; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_33_clock = clock;
  assign FP_multiplier_10ccs_33_reset = reset;
  assign FP_multiplier_10ccs_33_io_in_a = io_in_a_33; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_33_io_in_b = io_in_b_33; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_34_clock = clock;
  assign FP_multiplier_10ccs_34_reset = reset;
  assign FP_multiplier_10ccs_34_io_in_a = io_in_a_34; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_34_io_in_b = io_in_b_34; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_35_clock = clock;
  assign FP_multiplier_10ccs_35_reset = reset;
  assign FP_multiplier_10ccs_35_io_in_a = io_in_a_35; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_35_io_in_b = io_in_b_35; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_36_clock = clock;
  assign FP_multiplier_10ccs_36_reset = reset;
  assign FP_multiplier_10ccs_36_io_in_a = io_in_a_36; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_36_io_in_b = io_in_b_36; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_37_clock = clock;
  assign FP_multiplier_10ccs_37_reset = reset;
  assign FP_multiplier_10ccs_37_io_in_a = io_in_a_37; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_37_io_in_b = io_in_b_37; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_38_clock = clock;
  assign FP_multiplier_10ccs_38_reset = reset;
  assign FP_multiplier_10ccs_38_io_in_a = io_in_a_38; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_38_io_in_b = io_in_b_38; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_39_clock = clock;
  assign FP_multiplier_10ccs_39_reset = reset;
  assign FP_multiplier_10ccs_39_io_in_a = io_in_a_39; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_39_io_in_b = io_in_b_39; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_40_clock = clock;
  assign FP_multiplier_10ccs_40_reset = reset;
  assign FP_multiplier_10ccs_40_io_in_a = io_in_a_40; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_40_io_in_b = io_in_b_40; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_41_clock = clock;
  assign FP_multiplier_10ccs_41_reset = reset;
  assign FP_multiplier_10ccs_41_io_in_a = io_in_a_41; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_41_io_in_b = io_in_b_41; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_42_clock = clock;
  assign FP_multiplier_10ccs_42_reset = reset;
  assign FP_multiplier_10ccs_42_io_in_a = io_in_a_42; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_42_io_in_b = io_in_b_42; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_43_clock = clock;
  assign FP_multiplier_10ccs_43_reset = reset;
  assign FP_multiplier_10ccs_43_io_in_a = io_in_a_43; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_43_io_in_b = io_in_b_43; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_44_clock = clock;
  assign FP_multiplier_10ccs_44_reset = reset;
  assign FP_multiplier_10ccs_44_io_in_a = io_in_a_44; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_44_io_in_b = io_in_b_44; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_45_clock = clock;
  assign FP_multiplier_10ccs_45_reset = reset;
  assign FP_multiplier_10ccs_45_io_in_a = io_in_a_45; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_45_io_in_b = io_in_b_45; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_46_clock = clock;
  assign FP_multiplier_10ccs_46_reset = reset;
  assign FP_multiplier_10ccs_46_io_in_a = io_in_a_46; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_46_io_in_b = io_in_b_46; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_47_clock = clock;
  assign FP_multiplier_10ccs_47_reset = reset;
  assign FP_multiplier_10ccs_47_io_in_a = io_in_a_47; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_47_io_in_b = io_in_b_47; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_48_clock = clock;
  assign FP_multiplier_10ccs_48_reset = reset;
  assign FP_multiplier_10ccs_48_io_in_a = io_in_a_48; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_48_io_in_b = io_in_b_48; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_49_clock = clock;
  assign FP_multiplier_10ccs_49_reset = reset;
  assign FP_multiplier_10ccs_49_io_in_a = io_in_a_49; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_49_io_in_b = io_in_b_49; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_50_clock = clock;
  assign FP_multiplier_10ccs_50_reset = reset;
  assign FP_multiplier_10ccs_50_io_in_a = io_in_a_50; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_50_io_in_b = io_in_b_50; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_51_clock = clock;
  assign FP_multiplier_10ccs_51_reset = reset;
  assign FP_multiplier_10ccs_51_io_in_a = io_in_a_51; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_51_io_in_b = io_in_b_51; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_52_clock = clock;
  assign FP_multiplier_10ccs_52_reset = reset;
  assign FP_multiplier_10ccs_52_io_in_a = io_in_a_52; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_52_io_in_b = io_in_b_52; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_53_clock = clock;
  assign FP_multiplier_10ccs_53_reset = reset;
  assign FP_multiplier_10ccs_53_io_in_a = io_in_a_53; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_53_io_in_b = io_in_b_53; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_54_clock = clock;
  assign FP_multiplier_10ccs_54_reset = reset;
  assign FP_multiplier_10ccs_54_io_in_a = io_in_a_54; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_54_io_in_b = io_in_b_54; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_55_clock = clock;
  assign FP_multiplier_10ccs_55_reset = reset;
  assign FP_multiplier_10ccs_55_io_in_a = io_in_a_55; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_55_io_in_b = io_in_b_55; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_56_clock = clock;
  assign FP_multiplier_10ccs_56_reset = reset;
  assign FP_multiplier_10ccs_56_io_in_a = io_in_a_56; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_56_io_in_b = io_in_b_56; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_57_clock = clock;
  assign FP_multiplier_10ccs_57_reset = reset;
  assign FP_multiplier_10ccs_57_io_in_a = io_in_a_57; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_57_io_in_b = io_in_b_57; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_58_clock = clock;
  assign FP_multiplier_10ccs_58_reset = reset;
  assign FP_multiplier_10ccs_58_io_in_a = io_in_a_58; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_58_io_in_b = io_in_b_58; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_59_clock = clock;
  assign FP_multiplier_10ccs_59_reset = reset;
  assign FP_multiplier_10ccs_59_io_in_a = io_in_a_59; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_59_io_in_b = io_in_b_59; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_60_clock = clock;
  assign FP_multiplier_10ccs_60_reset = reset;
  assign FP_multiplier_10ccs_60_io_in_a = io_in_a_60; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_60_io_in_b = io_in_b_60; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_61_clock = clock;
  assign FP_multiplier_10ccs_61_reset = reset;
  assign FP_multiplier_10ccs_61_io_in_a = io_in_a_61; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_61_io_in_b = io_in_b_61; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_62_clock = clock;
  assign FP_multiplier_10ccs_62_reset = reset;
  assign FP_multiplier_10ccs_62_io_in_a = io_in_a_62; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_62_io_in_b = io_in_b_62; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_63_clock = clock;
  assign FP_multiplier_10ccs_63_reset = reset;
  assign FP_multiplier_10ccs_63_io_in_a = io_in_a_63; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_63_io_in_b = io_in_b_63; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_64_clock = clock;
  assign FP_multiplier_10ccs_64_reset = reset;
  assign FP_multiplier_10ccs_64_io_in_a = io_in_a_64; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_64_io_in_b = io_in_b_64; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_65_clock = clock;
  assign FP_multiplier_10ccs_65_reset = reset;
  assign FP_multiplier_10ccs_65_io_in_a = io_in_a_65; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_65_io_in_b = io_in_b_65; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_66_clock = clock;
  assign FP_multiplier_10ccs_66_reset = reset;
  assign FP_multiplier_10ccs_66_io_in_a = io_in_a_66; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_66_io_in_b = io_in_b_66; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_67_clock = clock;
  assign FP_multiplier_10ccs_67_reset = reset;
  assign FP_multiplier_10ccs_67_io_in_a = io_in_a_67; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_67_io_in_b = io_in_b_67; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_68_clock = clock;
  assign FP_multiplier_10ccs_68_reset = reset;
  assign FP_multiplier_10ccs_68_io_in_a = io_in_a_68; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_68_io_in_b = io_in_b_68; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_69_clock = clock;
  assign FP_multiplier_10ccs_69_reset = reset;
  assign FP_multiplier_10ccs_69_io_in_a = io_in_a_69; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_69_io_in_b = io_in_b_69; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_70_clock = clock;
  assign FP_multiplier_10ccs_70_reset = reset;
  assign FP_multiplier_10ccs_70_io_in_a = io_in_a_70; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_70_io_in_b = io_in_b_70; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_71_clock = clock;
  assign FP_multiplier_10ccs_71_reset = reset;
  assign FP_multiplier_10ccs_71_io_in_a = io_in_a_71; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_71_io_in_b = io_in_b_71; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_72_clock = clock;
  assign FP_multiplier_10ccs_72_reset = reset;
  assign FP_multiplier_10ccs_72_io_in_a = io_in_a_72; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_72_io_in_b = io_in_b_72; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_73_clock = clock;
  assign FP_multiplier_10ccs_73_reset = reset;
  assign FP_multiplier_10ccs_73_io_in_a = io_in_a_73; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_73_io_in_b = io_in_b_73; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_74_clock = clock;
  assign FP_multiplier_10ccs_74_reset = reset;
  assign FP_multiplier_10ccs_74_io_in_a = io_in_a_74; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_74_io_in_b = io_in_b_74; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_75_clock = clock;
  assign FP_multiplier_10ccs_75_reset = reset;
  assign FP_multiplier_10ccs_75_io_in_a = io_in_a_75; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_75_io_in_b = io_in_b_75; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_76_clock = clock;
  assign FP_multiplier_10ccs_76_reset = reset;
  assign FP_multiplier_10ccs_76_io_in_a = io_in_a_76; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_76_io_in_b = io_in_b_76; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_77_clock = clock;
  assign FP_multiplier_10ccs_77_reset = reset;
  assign FP_multiplier_10ccs_77_io_in_a = io_in_a_77; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_77_io_in_b = io_in_b_77; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_78_clock = clock;
  assign FP_multiplier_10ccs_78_reset = reset;
  assign FP_multiplier_10ccs_78_io_in_a = io_in_a_78; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_78_io_in_b = io_in_b_78; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_79_clock = clock;
  assign FP_multiplier_10ccs_79_reset = reset;
  assign FP_multiplier_10ccs_79_io_in_a = io_in_a_79; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_79_io_in_b = io_in_b_79; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_80_clock = clock;
  assign FP_multiplier_10ccs_80_reset = reset;
  assign FP_multiplier_10ccs_80_io_in_a = io_in_a_80; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_80_io_in_b = io_in_b_80; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_81_clock = clock;
  assign FP_multiplier_10ccs_81_reset = reset;
  assign FP_multiplier_10ccs_81_io_in_a = io_in_a_81; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_81_io_in_b = io_in_b_81; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_82_clock = clock;
  assign FP_multiplier_10ccs_82_reset = reset;
  assign FP_multiplier_10ccs_82_io_in_a = io_in_a_82; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_82_io_in_b = io_in_b_82; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_83_clock = clock;
  assign FP_multiplier_10ccs_83_reset = reset;
  assign FP_multiplier_10ccs_83_io_in_a = io_in_a_83; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_83_io_in_b = io_in_b_83; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_84_clock = clock;
  assign FP_multiplier_10ccs_84_reset = reset;
  assign FP_multiplier_10ccs_84_io_in_a = io_in_a_84; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_84_io_in_b = io_in_b_84; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_85_clock = clock;
  assign FP_multiplier_10ccs_85_reset = reset;
  assign FP_multiplier_10ccs_85_io_in_a = io_in_a_85; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_85_io_in_b = io_in_b_85; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_86_clock = clock;
  assign FP_multiplier_10ccs_86_reset = reset;
  assign FP_multiplier_10ccs_86_io_in_a = io_in_a_86; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_86_io_in_b = io_in_b_86; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_87_clock = clock;
  assign FP_multiplier_10ccs_87_reset = reset;
  assign FP_multiplier_10ccs_87_io_in_a = io_in_a_87; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_87_io_in_b = io_in_b_87; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_88_clock = clock;
  assign FP_multiplier_10ccs_88_reset = reset;
  assign FP_multiplier_10ccs_88_io_in_a = io_in_a_88; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_88_io_in_b = io_in_b_88; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_89_clock = clock;
  assign FP_multiplier_10ccs_89_reset = reset;
  assign FP_multiplier_10ccs_89_io_in_a = io_in_a_89; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_89_io_in_b = io_in_b_89; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_90_clock = clock;
  assign FP_multiplier_10ccs_90_reset = reset;
  assign FP_multiplier_10ccs_90_io_in_a = io_in_a_90; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_90_io_in_b = io_in_b_90; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_91_clock = clock;
  assign FP_multiplier_10ccs_91_reset = reset;
  assign FP_multiplier_10ccs_91_io_in_a = io_in_a_91; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_91_io_in_b = io_in_b_91; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_92_clock = clock;
  assign FP_multiplier_10ccs_92_reset = reset;
  assign FP_multiplier_10ccs_92_io_in_a = io_in_a_92; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_92_io_in_b = io_in_b_92; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_93_clock = clock;
  assign FP_multiplier_10ccs_93_reset = reset;
  assign FP_multiplier_10ccs_93_io_in_a = io_in_a_93; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_93_io_in_b = io_in_b_93; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_94_clock = clock;
  assign FP_multiplier_10ccs_94_reset = reset;
  assign FP_multiplier_10ccs_94_io_in_a = io_in_a_94; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_94_io_in_b = io_in_b_94; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_95_clock = clock;
  assign FP_multiplier_10ccs_95_reset = reset;
  assign FP_multiplier_10ccs_95_io_in_a = io_in_a_95; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_95_io_in_b = io_in_b_95; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_96_clock = clock;
  assign FP_multiplier_10ccs_96_reset = reset;
  assign FP_multiplier_10ccs_96_io_in_a = io_in_a_96; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_96_io_in_b = io_in_b_96; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_97_clock = clock;
  assign FP_multiplier_10ccs_97_reset = reset;
  assign FP_multiplier_10ccs_97_io_in_a = io_in_a_97; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_97_io_in_b = io_in_b_97; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_98_clock = clock;
  assign FP_multiplier_10ccs_98_reset = reset;
  assign FP_multiplier_10ccs_98_io_in_a = io_in_a_98; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_98_io_in_b = io_in_b_98; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_99_clock = clock;
  assign FP_multiplier_10ccs_99_reset = reset;
  assign FP_multiplier_10ccs_99_io_in_a = io_in_a_99; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_99_io_in_b = io_in_b_99; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_100_clock = clock;
  assign FP_multiplier_10ccs_100_reset = reset;
  assign FP_multiplier_10ccs_100_io_in_a = io_in_a_100; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_100_io_in_b = io_in_b_100; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_101_clock = clock;
  assign FP_multiplier_10ccs_101_reset = reset;
  assign FP_multiplier_10ccs_101_io_in_a = io_in_a_101; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_101_io_in_b = io_in_b_101; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_102_clock = clock;
  assign FP_multiplier_10ccs_102_reset = reset;
  assign FP_multiplier_10ccs_102_io_in_a = io_in_a_102; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_102_io_in_b = io_in_b_102; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_103_clock = clock;
  assign FP_multiplier_10ccs_103_reset = reset;
  assign FP_multiplier_10ccs_103_io_in_a = io_in_a_103; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_103_io_in_b = io_in_b_103; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_104_clock = clock;
  assign FP_multiplier_10ccs_104_reset = reset;
  assign FP_multiplier_10ccs_104_io_in_a = io_in_a_104; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_104_io_in_b = io_in_b_104; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_105_clock = clock;
  assign FP_multiplier_10ccs_105_reset = reset;
  assign FP_multiplier_10ccs_105_io_in_a = io_in_a_105; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_105_io_in_b = io_in_b_105; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_106_clock = clock;
  assign FP_multiplier_10ccs_106_reset = reset;
  assign FP_multiplier_10ccs_106_io_in_a = io_in_a_106; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_106_io_in_b = io_in_b_106; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_107_clock = clock;
  assign FP_multiplier_10ccs_107_reset = reset;
  assign FP_multiplier_10ccs_107_io_in_a = io_in_a_107; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_107_io_in_b = io_in_b_107; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_108_clock = clock;
  assign FP_multiplier_10ccs_108_reset = reset;
  assign FP_multiplier_10ccs_108_io_in_a = io_in_a_108; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_108_io_in_b = io_in_b_108; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_109_clock = clock;
  assign FP_multiplier_10ccs_109_reset = reset;
  assign FP_multiplier_10ccs_109_io_in_a = io_in_a_109; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_109_io_in_b = io_in_b_109; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_110_clock = clock;
  assign FP_multiplier_10ccs_110_reset = reset;
  assign FP_multiplier_10ccs_110_io_in_a = io_in_a_110; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_110_io_in_b = io_in_b_110; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_111_clock = clock;
  assign FP_multiplier_10ccs_111_reset = reset;
  assign FP_multiplier_10ccs_111_io_in_a = io_in_a_111; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_111_io_in_b = io_in_b_111; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_112_clock = clock;
  assign FP_multiplier_10ccs_112_reset = reset;
  assign FP_multiplier_10ccs_112_io_in_a = io_in_a_112; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_112_io_in_b = io_in_b_112; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_113_clock = clock;
  assign FP_multiplier_10ccs_113_reset = reset;
  assign FP_multiplier_10ccs_113_io_in_a = io_in_a_113; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_113_io_in_b = io_in_b_113; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_114_clock = clock;
  assign FP_multiplier_10ccs_114_reset = reset;
  assign FP_multiplier_10ccs_114_io_in_a = io_in_a_114; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_114_io_in_b = io_in_b_114; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_115_clock = clock;
  assign FP_multiplier_10ccs_115_reset = reset;
  assign FP_multiplier_10ccs_115_io_in_a = io_in_a_115; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_115_io_in_b = io_in_b_115; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_116_clock = clock;
  assign FP_multiplier_10ccs_116_reset = reset;
  assign FP_multiplier_10ccs_116_io_in_a = io_in_a_116; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_116_io_in_b = io_in_b_116; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_117_clock = clock;
  assign FP_multiplier_10ccs_117_reset = reset;
  assign FP_multiplier_10ccs_117_io_in_a = io_in_a_117; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_117_io_in_b = io_in_b_117; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_118_clock = clock;
  assign FP_multiplier_10ccs_118_reset = reset;
  assign FP_multiplier_10ccs_118_io_in_a = io_in_a_118; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_118_io_in_b = io_in_b_118; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_119_clock = clock;
  assign FP_multiplier_10ccs_119_reset = reset;
  assign FP_multiplier_10ccs_119_io_in_a = io_in_a_119; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_119_io_in_b = io_in_b_119; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_120_clock = clock;
  assign FP_multiplier_10ccs_120_reset = reset;
  assign FP_multiplier_10ccs_120_io_in_a = io_in_a_120; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_120_io_in_b = io_in_b_120; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_121_clock = clock;
  assign FP_multiplier_10ccs_121_reset = reset;
  assign FP_multiplier_10ccs_121_io_in_a = io_in_a_121; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_121_io_in_b = io_in_b_121; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_122_clock = clock;
  assign FP_multiplier_10ccs_122_reset = reset;
  assign FP_multiplier_10ccs_122_io_in_a = io_in_a_122; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_122_io_in_b = io_in_b_122; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_123_clock = clock;
  assign FP_multiplier_10ccs_123_reset = reset;
  assign FP_multiplier_10ccs_123_io_in_a = io_in_a_123; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_123_io_in_b = io_in_b_123; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_124_clock = clock;
  assign FP_multiplier_10ccs_124_reset = reset;
  assign FP_multiplier_10ccs_124_io_in_a = io_in_a_124; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_124_io_in_b = io_in_b_124; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_125_clock = clock;
  assign FP_multiplier_10ccs_125_reset = reset;
  assign FP_multiplier_10ccs_125_io_in_a = io_in_a_125; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_125_io_in_b = io_in_b_125; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_126_clock = clock;
  assign FP_multiplier_10ccs_126_reset = reset;
  assign FP_multiplier_10ccs_126_io_in_a = io_in_a_126; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_126_io_in_b = io_in_b_126; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_multiplier_10ccs_127_clock = clock;
  assign FP_multiplier_10ccs_127_reset = reset;
  assign FP_multiplier_10ccs_127_io_in_a = io_in_a_127; // @[FloatingPointDesigns.scala 2411:47]
  assign FP_multiplier_10ccs_127_io_in_b = io_in_b_127; // @[FloatingPointDesigns.scala 2412:47]
  assign FP_adder_13ccs_clock = clock;
  assign FP_adder_13ccs_reset = reset;
  assign FP_adder_13ccs_io_in_a = FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_io_in_b = FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_1_clock = clock;
  assign FP_adder_13ccs_1_reset = reset;
  assign FP_adder_13ccs_1_io_in_a = FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_1_io_in_b = FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_2_clock = clock;
  assign FP_adder_13ccs_2_reset = reset;
  assign FP_adder_13ccs_2_io_in_a = FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_2_io_in_b = FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_3_clock = clock;
  assign FP_adder_13ccs_3_reset = reset;
  assign FP_adder_13ccs_3_io_in_a = FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_3_io_in_b = FP_multiplier_10ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_4_clock = clock;
  assign FP_adder_13ccs_4_reset = reset;
  assign FP_adder_13ccs_4_io_in_a = FP_multiplier_10ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_4_io_in_b = FP_multiplier_10ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_5_clock = clock;
  assign FP_adder_13ccs_5_reset = reset;
  assign FP_adder_13ccs_5_io_in_a = FP_multiplier_10ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_5_io_in_b = FP_multiplier_10ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_6_clock = clock;
  assign FP_adder_13ccs_6_reset = reset;
  assign FP_adder_13ccs_6_io_in_a = FP_multiplier_10ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_6_io_in_b = FP_multiplier_10ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_7_clock = clock;
  assign FP_adder_13ccs_7_reset = reset;
  assign FP_adder_13ccs_7_io_in_a = FP_multiplier_10ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_7_io_in_b = FP_multiplier_10ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_8_clock = clock;
  assign FP_adder_13ccs_8_reset = reset;
  assign FP_adder_13ccs_8_io_in_a = FP_multiplier_10ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_8_io_in_b = FP_multiplier_10ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_9_clock = clock;
  assign FP_adder_13ccs_9_reset = reset;
  assign FP_adder_13ccs_9_io_in_a = FP_multiplier_10ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_9_io_in_b = FP_multiplier_10ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_10_clock = clock;
  assign FP_adder_13ccs_10_reset = reset;
  assign FP_adder_13ccs_10_io_in_a = FP_multiplier_10ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_10_io_in_b = FP_multiplier_10ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_11_clock = clock;
  assign FP_adder_13ccs_11_reset = reset;
  assign FP_adder_13ccs_11_io_in_a = FP_multiplier_10ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_11_io_in_b = FP_multiplier_10ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_12_clock = clock;
  assign FP_adder_13ccs_12_reset = reset;
  assign FP_adder_13ccs_12_io_in_a = FP_multiplier_10ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_12_io_in_b = FP_multiplier_10ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_13_clock = clock;
  assign FP_adder_13ccs_13_reset = reset;
  assign FP_adder_13ccs_13_io_in_a = FP_multiplier_10ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_13_io_in_b = FP_multiplier_10ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_14_clock = clock;
  assign FP_adder_13ccs_14_reset = reset;
  assign FP_adder_13ccs_14_io_in_a = FP_multiplier_10ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_14_io_in_b = FP_multiplier_10ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_15_clock = clock;
  assign FP_adder_13ccs_15_reset = reset;
  assign FP_adder_13ccs_15_io_in_a = FP_multiplier_10ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_15_io_in_b = FP_multiplier_10ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_16_clock = clock;
  assign FP_adder_13ccs_16_reset = reset;
  assign FP_adder_13ccs_16_io_in_a = FP_multiplier_10ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_16_io_in_b = FP_multiplier_10ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_17_clock = clock;
  assign FP_adder_13ccs_17_reset = reset;
  assign FP_adder_13ccs_17_io_in_a = FP_multiplier_10ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_17_io_in_b = FP_multiplier_10ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_18_clock = clock;
  assign FP_adder_13ccs_18_reset = reset;
  assign FP_adder_13ccs_18_io_in_a = FP_multiplier_10ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_18_io_in_b = FP_multiplier_10ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_19_clock = clock;
  assign FP_adder_13ccs_19_reset = reset;
  assign FP_adder_13ccs_19_io_in_a = FP_multiplier_10ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_19_io_in_b = FP_multiplier_10ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_20_clock = clock;
  assign FP_adder_13ccs_20_reset = reset;
  assign FP_adder_13ccs_20_io_in_a = FP_multiplier_10ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_20_io_in_b = FP_multiplier_10ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_21_clock = clock;
  assign FP_adder_13ccs_21_reset = reset;
  assign FP_adder_13ccs_21_io_in_a = FP_multiplier_10ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_21_io_in_b = FP_multiplier_10ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_22_clock = clock;
  assign FP_adder_13ccs_22_reset = reset;
  assign FP_adder_13ccs_22_io_in_a = FP_multiplier_10ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_22_io_in_b = FP_multiplier_10ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_23_clock = clock;
  assign FP_adder_13ccs_23_reset = reset;
  assign FP_adder_13ccs_23_io_in_a = FP_multiplier_10ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_23_io_in_b = FP_multiplier_10ccs_47_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_24_clock = clock;
  assign FP_adder_13ccs_24_reset = reset;
  assign FP_adder_13ccs_24_io_in_a = FP_multiplier_10ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_24_io_in_b = FP_multiplier_10ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_25_clock = clock;
  assign FP_adder_13ccs_25_reset = reset;
  assign FP_adder_13ccs_25_io_in_a = FP_multiplier_10ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_25_io_in_b = FP_multiplier_10ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_26_clock = clock;
  assign FP_adder_13ccs_26_reset = reset;
  assign FP_adder_13ccs_26_io_in_a = FP_multiplier_10ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_26_io_in_b = FP_multiplier_10ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_27_clock = clock;
  assign FP_adder_13ccs_27_reset = reset;
  assign FP_adder_13ccs_27_io_in_a = FP_multiplier_10ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_27_io_in_b = FP_multiplier_10ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_28_clock = clock;
  assign FP_adder_13ccs_28_reset = reset;
  assign FP_adder_13ccs_28_io_in_a = FP_multiplier_10ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_28_io_in_b = FP_multiplier_10ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_29_clock = clock;
  assign FP_adder_13ccs_29_reset = reset;
  assign FP_adder_13ccs_29_io_in_a = FP_multiplier_10ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_29_io_in_b = FP_multiplier_10ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_30_clock = clock;
  assign FP_adder_13ccs_30_reset = reset;
  assign FP_adder_13ccs_30_io_in_a = FP_multiplier_10ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_30_io_in_b = FP_multiplier_10ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_31_clock = clock;
  assign FP_adder_13ccs_31_reset = reset;
  assign FP_adder_13ccs_31_io_in_a = FP_multiplier_10ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_31_io_in_b = FP_multiplier_10ccs_63_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_32_clock = clock;
  assign FP_adder_13ccs_32_reset = reset;
  assign FP_adder_13ccs_32_io_in_a = FP_multiplier_10ccs_64_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_32_io_in_b = FP_multiplier_10ccs_65_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_33_clock = clock;
  assign FP_adder_13ccs_33_reset = reset;
  assign FP_adder_13ccs_33_io_in_a = FP_multiplier_10ccs_66_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_33_io_in_b = FP_multiplier_10ccs_67_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_34_clock = clock;
  assign FP_adder_13ccs_34_reset = reset;
  assign FP_adder_13ccs_34_io_in_a = FP_multiplier_10ccs_68_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_34_io_in_b = FP_multiplier_10ccs_69_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_35_clock = clock;
  assign FP_adder_13ccs_35_reset = reset;
  assign FP_adder_13ccs_35_io_in_a = FP_multiplier_10ccs_70_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_35_io_in_b = FP_multiplier_10ccs_71_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_36_clock = clock;
  assign FP_adder_13ccs_36_reset = reset;
  assign FP_adder_13ccs_36_io_in_a = FP_multiplier_10ccs_72_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_36_io_in_b = FP_multiplier_10ccs_73_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_37_clock = clock;
  assign FP_adder_13ccs_37_reset = reset;
  assign FP_adder_13ccs_37_io_in_a = FP_multiplier_10ccs_74_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_37_io_in_b = FP_multiplier_10ccs_75_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_38_clock = clock;
  assign FP_adder_13ccs_38_reset = reset;
  assign FP_adder_13ccs_38_io_in_a = FP_multiplier_10ccs_76_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_38_io_in_b = FP_multiplier_10ccs_77_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_39_clock = clock;
  assign FP_adder_13ccs_39_reset = reset;
  assign FP_adder_13ccs_39_io_in_a = FP_multiplier_10ccs_78_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_39_io_in_b = FP_multiplier_10ccs_79_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_40_clock = clock;
  assign FP_adder_13ccs_40_reset = reset;
  assign FP_adder_13ccs_40_io_in_a = FP_multiplier_10ccs_80_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_40_io_in_b = FP_multiplier_10ccs_81_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_41_clock = clock;
  assign FP_adder_13ccs_41_reset = reset;
  assign FP_adder_13ccs_41_io_in_a = FP_multiplier_10ccs_82_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_41_io_in_b = FP_multiplier_10ccs_83_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_42_clock = clock;
  assign FP_adder_13ccs_42_reset = reset;
  assign FP_adder_13ccs_42_io_in_a = FP_multiplier_10ccs_84_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_42_io_in_b = FP_multiplier_10ccs_85_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_43_clock = clock;
  assign FP_adder_13ccs_43_reset = reset;
  assign FP_adder_13ccs_43_io_in_a = FP_multiplier_10ccs_86_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_43_io_in_b = FP_multiplier_10ccs_87_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_44_clock = clock;
  assign FP_adder_13ccs_44_reset = reset;
  assign FP_adder_13ccs_44_io_in_a = FP_multiplier_10ccs_88_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_44_io_in_b = FP_multiplier_10ccs_89_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_45_clock = clock;
  assign FP_adder_13ccs_45_reset = reset;
  assign FP_adder_13ccs_45_io_in_a = FP_multiplier_10ccs_90_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_45_io_in_b = FP_multiplier_10ccs_91_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_46_clock = clock;
  assign FP_adder_13ccs_46_reset = reset;
  assign FP_adder_13ccs_46_io_in_a = FP_multiplier_10ccs_92_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_46_io_in_b = FP_multiplier_10ccs_93_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_47_clock = clock;
  assign FP_adder_13ccs_47_reset = reset;
  assign FP_adder_13ccs_47_io_in_a = FP_multiplier_10ccs_94_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_47_io_in_b = FP_multiplier_10ccs_95_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_48_clock = clock;
  assign FP_adder_13ccs_48_reset = reset;
  assign FP_adder_13ccs_48_io_in_a = FP_multiplier_10ccs_96_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_48_io_in_b = FP_multiplier_10ccs_97_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_49_clock = clock;
  assign FP_adder_13ccs_49_reset = reset;
  assign FP_adder_13ccs_49_io_in_a = FP_multiplier_10ccs_98_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_49_io_in_b = FP_multiplier_10ccs_99_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_50_clock = clock;
  assign FP_adder_13ccs_50_reset = reset;
  assign FP_adder_13ccs_50_io_in_a = FP_multiplier_10ccs_100_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_50_io_in_b = FP_multiplier_10ccs_101_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_51_clock = clock;
  assign FP_adder_13ccs_51_reset = reset;
  assign FP_adder_13ccs_51_io_in_a = FP_multiplier_10ccs_102_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_51_io_in_b = FP_multiplier_10ccs_103_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_52_clock = clock;
  assign FP_adder_13ccs_52_reset = reset;
  assign FP_adder_13ccs_52_io_in_a = FP_multiplier_10ccs_104_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_52_io_in_b = FP_multiplier_10ccs_105_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_53_clock = clock;
  assign FP_adder_13ccs_53_reset = reset;
  assign FP_adder_13ccs_53_io_in_a = FP_multiplier_10ccs_106_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_53_io_in_b = FP_multiplier_10ccs_107_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_54_clock = clock;
  assign FP_adder_13ccs_54_reset = reset;
  assign FP_adder_13ccs_54_io_in_a = FP_multiplier_10ccs_108_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_54_io_in_b = FP_multiplier_10ccs_109_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_55_clock = clock;
  assign FP_adder_13ccs_55_reset = reset;
  assign FP_adder_13ccs_55_io_in_a = FP_multiplier_10ccs_110_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_55_io_in_b = FP_multiplier_10ccs_111_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_56_clock = clock;
  assign FP_adder_13ccs_56_reset = reset;
  assign FP_adder_13ccs_56_io_in_a = FP_multiplier_10ccs_112_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_56_io_in_b = FP_multiplier_10ccs_113_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_57_clock = clock;
  assign FP_adder_13ccs_57_reset = reset;
  assign FP_adder_13ccs_57_io_in_a = FP_multiplier_10ccs_114_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_57_io_in_b = FP_multiplier_10ccs_115_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_58_clock = clock;
  assign FP_adder_13ccs_58_reset = reset;
  assign FP_adder_13ccs_58_io_in_a = FP_multiplier_10ccs_116_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_58_io_in_b = FP_multiplier_10ccs_117_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_59_clock = clock;
  assign FP_adder_13ccs_59_reset = reset;
  assign FP_adder_13ccs_59_io_in_a = FP_multiplier_10ccs_118_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_59_io_in_b = FP_multiplier_10ccs_119_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_60_clock = clock;
  assign FP_adder_13ccs_60_reset = reset;
  assign FP_adder_13ccs_60_io_in_a = FP_multiplier_10ccs_120_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_60_io_in_b = FP_multiplier_10ccs_121_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_61_clock = clock;
  assign FP_adder_13ccs_61_reset = reset;
  assign FP_adder_13ccs_61_io_in_a = FP_multiplier_10ccs_122_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_61_io_in_b = FP_multiplier_10ccs_123_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_62_clock = clock;
  assign FP_adder_13ccs_62_reset = reset;
  assign FP_adder_13ccs_62_io_in_a = FP_multiplier_10ccs_124_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_62_io_in_b = FP_multiplier_10ccs_125_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_63_clock = clock;
  assign FP_adder_13ccs_63_reset = reset;
  assign FP_adder_13ccs_63_io_in_a = FP_multiplier_10ccs_126_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_63_io_in_b = FP_multiplier_10ccs_127_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_64_clock = clock;
  assign FP_adder_13ccs_64_reset = reset;
  assign FP_adder_13ccs_64_io_in_a = FP_adder_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_64_io_in_b = FP_adder_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_65_clock = clock;
  assign FP_adder_13ccs_65_reset = reset;
  assign FP_adder_13ccs_65_io_in_a = FP_adder_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_65_io_in_b = FP_adder_13ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_66_clock = clock;
  assign FP_adder_13ccs_66_reset = reset;
  assign FP_adder_13ccs_66_io_in_a = FP_adder_13ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_66_io_in_b = FP_adder_13ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_67_clock = clock;
  assign FP_adder_13ccs_67_reset = reset;
  assign FP_adder_13ccs_67_io_in_a = FP_adder_13ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_67_io_in_b = FP_adder_13ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_68_clock = clock;
  assign FP_adder_13ccs_68_reset = reset;
  assign FP_adder_13ccs_68_io_in_a = FP_adder_13ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_68_io_in_b = FP_adder_13ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_69_clock = clock;
  assign FP_adder_13ccs_69_reset = reset;
  assign FP_adder_13ccs_69_io_in_a = FP_adder_13ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_69_io_in_b = FP_adder_13ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_70_clock = clock;
  assign FP_adder_13ccs_70_reset = reset;
  assign FP_adder_13ccs_70_io_in_a = FP_adder_13ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_70_io_in_b = FP_adder_13ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_71_clock = clock;
  assign FP_adder_13ccs_71_reset = reset;
  assign FP_adder_13ccs_71_io_in_a = FP_adder_13ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_71_io_in_b = FP_adder_13ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_72_clock = clock;
  assign FP_adder_13ccs_72_reset = reset;
  assign FP_adder_13ccs_72_io_in_a = FP_adder_13ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_72_io_in_b = FP_adder_13ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_73_clock = clock;
  assign FP_adder_13ccs_73_reset = reset;
  assign FP_adder_13ccs_73_io_in_a = FP_adder_13ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_73_io_in_b = FP_adder_13ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_74_clock = clock;
  assign FP_adder_13ccs_74_reset = reset;
  assign FP_adder_13ccs_74_io_in_a = FP_adder_13ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_74_io_in_b = FP_adder_13ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_75_clock = clock;
  assign FP_adder_13ccs_75_reset = reset;
  assign FP_adder_13ccs_75_io_in_a = FP_adder_13ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_75_io_in_b = FP_adder_13ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_76_clock = clock;
  assign FP_adder_13ccs_76_reset = reset;
  assign FP_adder_13ccs_76_io_in_a = FP_adder_13ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_76_io_in_b = FP_adder_13ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_77_clock = clock;
  assign FP_adder_13ccs_77_reset = reset;
  assign FP_adder_13ccs_77_io_in_a = FP_adder_13ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_77_io_in_b = FP_adder_13ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_78_clock = clock;
  assign FP_adder_13ccs_78_reset = reset;
  assign FP_adder_13ccs_78_io_in_a = FP_adder_13ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_78_io_in_b = FP_adder_13ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_79_clock = clock;
  assign FP_adder_13ccs_79_reset = reset;
  assign FP_adder_13ccs_79_io_in_a = FP_adder_13ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_79_io_in_b = FP_adder_13ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_80_clock = clock;
  assign FP_adder_13ccs_80_reset = reset;
  assign FP_adder_13ccs_80_io_in_a = FP_adder_13ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_80_io_in_b = FP_adder_13ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_81_clock = clock;
  assign FP_adder_13ccs_81_reset = reset;
  assign FP_adder_13ccs_81_io_in_a = FP_adder_13ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_81_io_in_b = FP_adder_13ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_82_clock = clock;
  assign FP_adder_13ccs_82_reset = reset;
  assign FP_adder_13ccs_82_io_in_a = FP_adder_13ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_82_io_in_b = FP_adder_13ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_83_clock = clock;
  assign FP_adder_13ccs_83_reset = reset;
  assign FP_adder_13ccs_83_io_in_a = FP_adder_13ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_83_io_in_b = FP_adder_13ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_84_clock = clock;
  assign FP_adder_13ccs_84_reset = reset;
  assign FP_adder_13ccs_84_io_in_a = FP_adder_13ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_84_io_in_b = FP_adder_13ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_85_clock = clock;
  assign FP_adder_13ccs_85_reset = reset;
  assign FP_adder_13ccs_85_io_in_a = FP_adder_13ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_85_io_in_b = FP_adder_13ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_86_clock = clock;
  assign FP_adder_13ccs_86_reset = reset;
  assign FP_adder_13ccs_86_io_in_a = FP_adder_13ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_86_io_in_b = FP_adder_13ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_87_clock = clock;
  assign FP_adder_13ccs_87_reset = reset;
  assign FP_adder_13ccs_87_io_in_a = FP_adder_13ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_87_io_in_b = FP_adder_13ccs_47_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_88_clock = clock;
  assign FP_adder_13ccs_88_reset = reset;
  assign FP_adder_13ccs_88_io_in_a = FP_adder_13ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_88_io_in_b = FP_adder_13ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_89_clock = clock;
  assign FP_adder_13ccs_89_reset = reset;
  assign FP_adder_13ccs_89_io_in_a = FP_adder_13ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_89_io_in_b = FP_adder_13ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_90_clock = clock;
  assign FP_adder_13ccs_90_reset = reset;
  assign FP_adder_13ccs_90_io_in_a = FP_adder_13ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_90_io_in_b = FP_adder_13ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_91_clock = clock;
  assign FP_adder_13ccs_91_reset = reset;
  assign FP_adder_13ccs_91_io_in_a = FP_adder_13ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_91_io_in_b = FP_adder_13ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_92_clock = clock;
  assign FP_adder_13ccs_92_reset = reset;
  assign FP_adder_13ccs_92_io_in_a = FP_adder_13ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_92_io_in_b = FP_adder_13ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_93_clock = clock;
  assign FP_adder_13ccs_93_reset = reset;
  assign FP_adder_13ccs_93_io_in_a = FP_adder_13ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_93_io_in_b = FP_adder_13ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_94_clock = clock;
  assign FP_adder_13ccs_94_reset = reset;
  assign FP_adder_13ccs_94_io_in_a = FP_adder_13ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_94_io_in_b = FP_adder_13ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_95_clock = clock;
  assign FP_adder_13ccs_95_reset = reset;
  assign FP_adder_13ccs_95_io_in_a = FP_adder_13ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_95_io_in_b = FP_adder_13ccs_63_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_96_clock = clock;
  assign FP_adder_13ccs_96_reset = reset;
  assign FP_adder_13ccs_96_io_in_a = FP_adder_13ccs_64_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_96_io_in_b = FP_adder_13ccs_65_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_97_clock = clock;
  assign FP_adder_13ccs_97_reset = reset;
  assign FP_adder_13ccs_97_io_in_a = FP_adder_13ccs_66_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_97_io_in_b = FP_adder_13ccs_67_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_98_clock = clock;
  assign FP_adder_13ccs_98_reset = reset;
  assign FP_adder_13ccs_98_io_in_a = FP_adder_13ccs_68_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_98_io_in_b = FP_adder_13ccs_69_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_99_clock = clock;
  assign FP_adder_13ccs_99_reset = reset;
  assign FP_adder_13ccs_99_io_in_a = FP_adder_13ccs_70_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_99_io_in_b = FP_adder_13ccs_71_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_100_clock = clock;
  assign FP_adder_13ccs_100_reset = reset;
  assign FP_adder_13ccs_100_io_in_a = FP_adder_13ccs_72_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_100_io_in_b = FP_adder_13ccs_73_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_101_clock = clock;
  assign FP_adder_13ccs_101_reset = reset;
  assign FP_adder_13ccs_101_io_in_a = FP_adder_13ccs_74_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_101_io_in_b = FP_adder_13ccs_75_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_102_clock = clock;
  assign FP_adder_13ccs_102_reset = reset;
  assign FP_adder_13ccs_102_io_in_a = FP_adder_13ccs_76_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_102_io_in_b = FP_adder_13ccs_77_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_103_clock = clock;
  assign FP_adder_13ccs_103_reset = reset;
  assign FP_adder_13ccs_103_io_in_a = FP_adder_13ccs_78_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_103_io_in_b = FP_adder_13ccs_79_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_104_clock = clock;
  assign FP_adder_13ccs_104_reset = reset;
  assign FP_adder_13ccs_104_io_in_a = FP_adder_13ccs_80_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_104_io_in_b = FP_adder_13ccs_81_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_105_clock = clock;
  assign FP_adder_13ccs_105_reset = reset;
  assign FP_adder_13ccs_105_io_in_a = FP_adder_13ccs_82_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_105_io_in_b = FP_adder_13ccs_83_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_106_clock = clock;
  assign FP_adder_13ccs_106_reset = reset;
  assign FP_adder_13ccs_106_io_in_a = FP_adder_13ccs_84_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_106_io_in_b = FP_adder_13ccs_85_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_107_clock = clock;
  assign FP_adder_13ccs_107_reset = reset;
  assign FP_adder_13ccs_107_io_in_a = FP_adder_13ccs_86_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_107_io_in_b = FP_adder_13ccs_87_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_108_clock = clock;
  assign FP_adder_13ccs_108_reset = reset;
  assign FP_adder_13ccs_108_io_in_a = FP_adder_13ccs_88_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_108_io_in_b = FP_adder_13ccs_89_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_109_clock = clock;
  assign FP_adder_13ccs_109_reset = reset;
  assign FP_adder_13ccs_109_io_in_a = FP_adder_13ccs_90_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_109_io_in_b = FP_adder_13ccs_91_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_110_clock = clock;
  assign FP_adder_13ccs_110_reset = reset;
  assign FP_adder_13ccs_110_io_in_a = FP_adder_13ccs_92_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_110_io_in_b = FP_adder_13ccs_93_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_111_clock = clock;
  assign FP_adder_13ccs_111_reset = reset;
  assign FP_adder_13ccs_111_io_in_a = FP_adder_13ccs_94_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_111_io_in_b = FP_adder_13ccs_95_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_112_clock = clock;
  assign FP_adder_13ccs_112_reset = reset;
  assign FP_adder_13ccs_112_io_in_a = FP_adder_13ccs_96_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_112_io_in_b = FP_adder_13ccs_97_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_113_clock = clock;
  assign FP_adder_13ccs_113_reset = reset;
  assign FP_adder_13ccs_113_io_in_a = FP_adder_13ccs_98_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_113_io_in_b = FP_adder_13ccs_99_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_114_clock = clock;
  assign FP_adder_13ccs_114_reset = reset;
  assign FP_adder_13ccs_114_io_in_a = FP_adder_13ccs_100_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_114_io_in_b = FP_adder_13ccs_101_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_115_clock = clock;
  assign FP_adder_13ccs_115_reset = reset;
  assign FP_adder_13ccs_115_io_in_a = FP_adder_13ccs_102_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_115_io_in_b = FP_adder_13ccs_103_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_116_clock = clock;
  assign FP_adder_13ccs_116_reset = reset;
  assign FP_adder_13ccs_116_io_in_a = FP_adder_13ccs_104_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_116_io_in_b = FP_adder_13ccs_105_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_117_clock = clock;
  assign FP_adder_13ccs_117_reset = reset;
  assign FP_adder_13ccs_117_io_in_a = FP_adder_13ccs_106_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_117_io_in_b = FP_adder_13ccs_107_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_118_clock = clock;
  assign FP_adder_13ccs_118_reset = reset;
  assign FP_adder_13ccs_118_io_in_a = FP_adder_13ccs_108_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_118_io_in_b = FP_adder_13ccs_109_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_119_clock = clock;
  assign FP_adder_13ccs_119_reset = reset;
  assign FP_adder_13ccs_119_io_in_a = FP_adder_13ccs_110_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_119_io_in_b = FP_adder_13ccs_111_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_120_clock = clock;
  assign FP_adder_13ccs_120_reset = reset;
  assign FP_adder_13ccs_120_io_in_a = FP_adder_13ccs_112_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_120_io_in_b = FP_adder_13ccs_113_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_121_clock = clock;
  assign FP_adder_13ccs_121_reset = reset;
  assign FP_adder_13ccs_121_io_in_a = FP_adder_13ccs_114_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_121_io_in_b = FP_adder_13ccs_115_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_122_clock = clock;
  assign FP_adder_13ccs_122_reset = reset;
  assign FP_adder_13ccs_122_io_in_a = FP_adder_13ccs_116_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_122_io_in_b = FP_adder_13ccs_117_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_123_clock = clock;
  assign FP_adder_13ccs_123_reset = reset;
  assign FP_adder_13ccs_123_io_in_a = FP_adder_13ccs_118_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_123_io_in_b = FP_adder_13ccs_119_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_124_clock = clock;
  assign FP_adder_13ccs_124_reset = reset;
  assign FP_adder_13ccs_124_io_in_a = FP_adder_13ccs_120_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_124_io_in_b = FP_adder_13ccs_121_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_125_clock = clock;
  assign FP_adder_13ccs_125_reset = reset;
  assign FP_adder_13ccs_125_io_in_a = FP_adder_13ccs_122_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_125_io_in_b = FP_adder_13ccs_123_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
  assign FP_adder_13ccs_126_clock = clock;
  assign FP_adder_13ccs_126_reset = reset;
  assign FP_adder_13ccs_126_io_in_a = FP_adder_13ccs_124_io_out_s; // @[FloatingPointDesigns.scala 2448:43]
  assign FP_adder_13ccs_126_io_in_b = FP_adder_13ccs_125_io_out_s; // @[FloatingPointDesigns.scala 2449:43]
endmodule
module FP_subtractor_13ccs(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
  wire  FP_adder_clock; // @[FloatingPointDesigns.scala 1650:26]
  wire  FP_adder_reset; // @[FloatingPointDesigns.scala 1650:26]
  wire [31:0] FP_adder_io_in_a; // @[FloatingPointDesigns.scala 1650:26]
  wire [31:0] FP_adder_io_in_b; // @[FloatingPointDesigns.scala 1650:26]
  wire [31:0] FP_adder_io_out_s; // @[FloatingPointDesigns.scala 1650:26]
  wire  _adjusted_in_b_T_1 = ~io_in_b[31]; // @[FloatingPointDesigns.scala 1653:23]
  FP_adder_13ccs FP_adder ( // @[FloatingPointDesigns.scala 1650:26]
    .clock(FP_adder_clock),
    .reset(FP_adder_reset),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  assign io_out_s = FP_adder_io_out_s; // @[FloatingPointDesigns.scala 1657:14]
  assign FP_adder_clock = clock;
  assign FP_adder_reset = reset;
  assign FP_adder_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 1655:22]
  assign FP_adder_io_in_b = {_adjusted_in_b_T_1,io_in_b[30:0]}; // @[FloatingPointDesigns.scala 1653:41]
endmodule
module FP_square_root_newfpu(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
`endif // RANDOMIZE_REG_INIT
  wire  FP_multiplier_10ccs_clock; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_multiplier_10ccs_reset; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_io_in_a; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_io_in_b; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_multiplier_10ccs_1_clock; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_multiplier_10ccs_1_reset; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_1_io_in_a; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_1_io_in_b; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_multiplier_10ccs_2_clock; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_multiplier_10ccs_2_reset; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_2_io_in_a; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_2_io_in_b; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_multiplier_10ccs_3_clock; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_multiplier_10ccs_3_reset; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_3_io_in_a; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_3_io_in_b; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_multiplier_10ccs_4_clock; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_multiplier_10ccs_4_reset; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_4_io_in_a; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_4_io_in_b; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_multiplier_10ccs_5_clock; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_multiplier_10ccs_5_reset; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_5_io_in_a; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_5_io_in_b; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_multiplier_10ccs_6_clock; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_multiplier_10ccs_6_reset; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_6_io_in_a; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_6_io_in_b; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_multiplier_10ccs_7_clock; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_multiplier_10ccs_7_reset; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_7_io_in_a; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_7_io_in_b; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_7_io_out_s; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_multiplier_10ccs_8_clock; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_multiplier_10ccs_8_reset; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_8_io_in_a; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_8_io_in_b; // @[FloatingPointDesigns.scala 1876:65]
  wire [31:0] FP_multiplier_10ccs_8_io_out_s; // @[FloatingPointDesigns.scala 1876:65]
  wire  FP_subtractor_13ccs_clock; // @[FloatingPointDesigns.scala 1877:50]
  wire  FP_subtractor_13ccs_reset; // @[FloatingPointDesigns.scala 1877:50]
  wire [31:0] FP_subtractor_13ccs_io_in_a; // @[FloatingPointDesigns.scala 1877:50]
  wire [31:0] FP_subtractor_13ccs_io_in_b; // @[FloatingPointDesigns.scala 1877:50]
  wire [31:0] FP_subtractor_13ccs_io_out_s; // @[FloatingPointDesigns.scala 1877:50]
  wire  FP_subtractor_13ccs_1_clock; // @[FloatingPointDesigns.scala 1877:50]
  wire  FP_subtractor_13ccs_1_reset; // @[FloatingPointDesigns.scala 1877:50]
  wire [31:0] FP_subtractor_13ccs_1_io_in_a; // @[FloatingPointDesigns.scala 1877:50]
  wire [31:0] FP_subtractor_13ccs_1_io_in_b; // @[FloatingPointDesigns.scala 1877:50]
  wire [31:0] FP_subtractor_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 1877:50]
  wire  FP_subtractor_13ccs_2_clock; // @[FloatingPointDesigns.scala 1877:50]
  wire  FP_subtractor_13ccs_2_reset; // @[FloatingPointDesigns.scala 1877:50]
  wire [31:0] FP_subtractor_13ccs_2_io_in_a; // @[FloatingPointDesigns.scala 1877:50]
  wire [31:0] FP_subtractor_13ccs_2_io_in_b; // @[FloatingPointDesigns.scala 1877:50]
  wire [31:0] FP_subtractor_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 1877:50]
  wire  multiplier4_clock; // @[FloatingPointDesigns.scala 1945:29]
  wire  multiplier4_reset; // @[FloatingPointDesigns.scala 1945:29]
  wire [31:0] multiplier4_io_in_a; // @[FloatingPointDesigns.scala 1945:29]
  wire [31:0] multiplier4_io_in_b; // @[FloatingPointDesigns.scala 1945:29]
  wire [31:0] multiplier4_io_out_s; // @[FloatingPointDesigns.scala 1945:29]
  wire [30:0] _number_T_1 = {{1'd0}, io_in_a[30:1]}; // @[FloatingPointDesigns.scala 1860:36]
  wire [30:0] _GEN_0 = io_in_a[30:0] > 31'h7ef477d4 ? 31'h3f7a3bea : _number_T_1; // @[FloatingPointDesigns.scala 1857:46 1858:14 1860:14]
  wire [31:0] number = {{1'd0}, _GEN_0}; // @[FloatingPointDesigns.scala 1854:22]
  wire [31:0] result = 32'h5f3759df - number; // @[FloatingPointDesigns.scala 1867:25]
  reg [31:0] x_n_0; // @[FloatingPointDesigns.scala 1869:22]
  reg [31:0] x_n_1; // @[FloatingPointDesigns.scala 1869:22]
  reg [31:0] x_n_2; // @[FloatingPointDesigns.scala 1869:22]
  reg [31:0] x_n_4; // @[FloatingPointDesigns.scala 1869:22]
  reg [31:0] x_n_5; // @[FloatingPointDesigns.scala 1869:22]
  reg [31:0] x_n_6; // @[FloatingPointDesigns.scala 1869:22]
  reg [31:0] x_n_8; // @[FloatingPointDesigns.scala 1869:22]
  reg [31:0] x_n_9; // @[FloatingPointDesigns.scala 1869:22]
  reg [31:0] x_n_10; // @[FloatingPointDesigns.scala 1869:22]
  reg [31:0] a_2_0; // @[FloatingPointDesigns.scala 1870:22]
  reg [31:0] a_2_1; // @[FloatingPointDesigns.scala 1870:22]
  reg [31:0] a_2_2; // @[FloatingPointDesigns.scala 1870:22]
  reg [31:0] a_2_3; // @[FloatingPointDesigns.scala 1870:22]
  reg [31:0] a_2_4; // @[FloatingPointDesigns.scala 1870:22]
  reg [31:0] a_2_5; // @[FloatingPointDesigns.scala 1870:22]
  reg [31:0] a_2_6; // @[FloatingPointDesigns.scala 1870:22]
  reg [31:0] a_2_7; // @[FloatingPointDesigns.scala 1870:22]
  reg [31:0] a_2_8; // @[FloatingPointDesigns.scala 1870:22]
  reg [31:0] a_2_9; // @[FloatingPointDesigns.scala 1870:22]
  reg [31:0] a_2_10; // @[FloatingPointDesigns.scala 1870:22]
  reg [31:0] a_2_11; // @[FloatingPointDesigns.scala 1870:22]
  reg [31:0] stage1_regs_0_0_0; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_0_0_1; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_0_0_2; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_0_0_3; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_0_0_4; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_0_0_5; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_0_0_6; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_0_0_7; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_0_0_8; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_0_1_0; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_0_1_1; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_0_1_2; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_0_1_3; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_0_1_4; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_0_1_5; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_0_1_6; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_0_1_7; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_0_1_8; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_0_0; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_0_1; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_0_2; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_0_3; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_0_4; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_0_5; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_0_6; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_0_7; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_0_8; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_1_0; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_1_1; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_1_2; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_1_3; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_1_4; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_1_5; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_1_6; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_1_7; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_1_1_8; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_0_0; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_0_1; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_0_2; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_0_3; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_0_4; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_0_5; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_0_6; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_0_7; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_0_8; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_1_0; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_1_1; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_1_2; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_1_3; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_1_4; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_1_5; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_1_6; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_1_7; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage1_regs_2_1_8; // @[FloatingPointDesigns.scala 1871:30]
  reg [31:0] stage2_regs_0_0_0; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_0_0_1; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_0_0_2; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_0_0_3; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_0_0_4; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_0_0_5; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_0_0_6; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_0_0_7; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_0_0_8; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_0_1_0; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_0_1_1; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_0_1_2; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_0_1_3; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_0_1_4; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_0_1_5; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_0_1_6; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_0_1_7; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_0_1_8; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_0_0; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_0_1; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_0_2; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_0_3; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_0_4; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_0_5; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_0_6; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_0_7; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_0_8; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_1_0; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_1_1; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_1_2; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_1_3; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_1_4; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_1_5; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_1_6; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_1_7; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_1_1_8; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_0_0; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_0_1; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_0_2; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_0_3; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_0_4; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_0_5; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_0_6; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_0_7; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_0_8; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_1_0; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_1_1; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_1_2; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_1_3; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_1_4; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_1_5; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_1_6; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_1_7; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage2_regs_2_1_8; // @[FloatingPointDesigns.scala 1872:30]
  reg [31:0] stage3_regs_0_0_0; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_0_1; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_0_2; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_0_3; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_0_4; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_0_5; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_0_6; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_0_7; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_0_8; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_0_9; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_0_10; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_0_11; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_1_0; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_1_1; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_1_2; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_1_3; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_1_4; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_1_5; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_1_6; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_1_7; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_1_8; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_1_9; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_1_10; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_0_1_11; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_0_0; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_0_1; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_0_2; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_0_3; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_0_4; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_0_5; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_0_6; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_0_7; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_0_8; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_0_9; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_0_10; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_0_11; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_1_0; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_1_1; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_1_2; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_1_3; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_1_4; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_1_5; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_1_6; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_1_7; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_1_8; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_1_9; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_1_10; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_1_1_11; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_0_0; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_0_1; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_0_2; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_0_3; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_0_4; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_0_5; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_0_6; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_0_7; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_0_8; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_0_9; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_0_10; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_0_11; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_1_0; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_1_1; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_1_2; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_1_3; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_1_4; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_1_5; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_1_6; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_1_7; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_1_8; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_1_9; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_1_10; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage3_regs_2_1_11; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage4_regs_0_1_0; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_0_1_1; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_0_1_2; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_0_1_3; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_0_1_4; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_0_1_5; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_0_1_6; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_0_1_7; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_0_1_8; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_1_1_0; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_1_1_1; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_1_1_2; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_1_1_3; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_1_1_4; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_1_1_5; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_1_1_6; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_1_1_7; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_1_1_8; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_2_1_0; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_2_1_1; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_2_1_2; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_2_1_3; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_2_1_4; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_2_1_5; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_2_1_6; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_2_1_7; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage4_regs_2_1_8; // @[FloatingPointDesigns.scala 1874:30]
  wire [7:0] _a_2_0_T_3 = io_in_a[30:23] - 8'h1; // @[FloatingPointDesigns.scala 1899:75]
  wire [31:0] _a_2_0_T_6 = {io_in_a[31],_a_2_0_T_3,io_in_a[22:0]}; // @[FloatingPointDesigns.scala 1899:82]
  wire [31:0] _GEN_139 = FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 1869:22 1906:28 1907:26]
  wire [31:0] _GEN_215 = FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 1869:22 1906:28 1907:26]
  wire [7:0] _restore_a_T_3 = stage4_regs_2_1_8[30:23] + 8'h1; // @[FloatingPointDesigns.scala 1944:106]
  wire [8:0] _restore_a_T_4 = {stage4_regs_2_1_8[31],_restore_a_T_3}; // @[FloatingPointDesigns.scala 1944:55]
  FP_multiplier_10ccs FP_multiplier_10ccs ( // @[FloatingPointDesigns.scala 1876:65]
    .clock(FP_multiplier_10ccs_clock),
    .reset(FP_multiplier_10ccs_reset),
    .io_in_a(FP_multiplier_10ccs_io_in_a),
    .io_in_b(FP_multiplier_10ccs_io_in_b),
    .io_out_s(FP_multiplier_10ccs_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_1 ( // @[FloatingPointDesigns.scala 1876:65]
    .clock(FP_multiplier_10ccs_1_clock),
    .reset(FP_multiplier_10ccs_1_reset),
    .io_in_a(FP_multiplier_10ccs_1_io_in_a),
    .io_in_b(FP_multiplier_10ccs_1_io_in_b),
    .io_out_s(FP_multiplier_10ccs_1_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_2 ( // @[FloatingPointDesigns.scala 1876:65]
    .clock(FP_multiplier_10ccs_2_clock),
    .reset(FP_multiplier_10ccs_2_reset),
    .io_in_a(FP_multiplier_10ccs_2_io_in_a),
    .io_in_b(FP_multiplier_10ccs_2_io_in_b),
    .io_out_s(FP_multiplier_10ccs_2_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_3 ( // @[FloatingPointDesigns.scala 1876:65]
    .clock(FP_multiplier_10ccs_3_clock),
    .reset(FP_multiplier_10ccs_3_reset),
    .io_in_a(FP_multiplier_10ccs_3_io_in_a),
    .io_in_b(FP_multiplier_10ccs_3_io_in_b),
    .io_out_s(FP_multiplier_10ccs_3_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_4 ( // @[FloatingPointDesigns.scala 1876:65]
    .clock(FP_multiplier_10ccs_4_clock),
    .reset(FP_multiplier_10ccs_4_reset),
    .io_in_a(FP_multiplier_10ccs_4_io_in_a),
    .io_in_b(FP_multiplier_10ccs_4_io_in_b),
    .io_out_s(FP_multiplier_10ccs_4_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_5 ( // @[FloatingPointDesigns.scala 1876:65]
    .clock(FP_multiplier_10ccs_5_clock),
    .reset(FP_multiplier_10ccs_5_reset),
    .io_in_a(FP_multiplier_10ccs_5_io_in_a),
    .io_in_b(FP_multiplier_10ccs_5_io_in_b),
    .io_out_s(FP_multiplier_10ccs_5_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_6 ( // @[FloatingPointDesigns.scala 1876:65]
    .clock(FP_multiplier_10ccs_6_clock),
    .reset(FP_multiplier_10ccs_6_reset),
    .io_in_a(FP_multiplier_10ccs_6_io_in_a),
    .io_in_b(FP_multiplier_10ccs_6_io_in_b),
    .io_out_s(FP_multiplier_10ccs_6_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_7 ( // @[FloatingPointDesigns.scala 1876:65]
    .clock(FP_multiplier_10ccs_7_clock),
    .reset(FP_multiplier_10ccs_7_reset),
    .io_in_a(FP_multiplier_10ccs_7_io_in_a),
    .io_in_b(FP_multiplier_10ccs_7_io_in_b),
    .io_out_s(FP_multiplier_10ccs_7_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_8 ( // @[FloatingPointDesigns.scala 1876:65]
    .clock(FP_multiplier_10ccs_8_clock),
    .reset(FP_multiplier_10ccs_8_reset),
    .io_in_a(FP_multiplier_10ccs_8_io_in_a),
    .io_in_b(FP_multiplier_10ccs_8_io_in_b),
    .io_out_s(FP_multiplier_10ccs_8_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs ( // @[FloatingPointDesigns.scala 1877:50]
    .clock(FP_subtractor_13ccs_clock),
    .reset(FP_subtractor_13ccs_reset),
    .io_in_a(FP_subtractor_13ccs_io_in_a),
    .io_in_b(FP_subtractor_13ccs_io_in_b),
    .io_out_s(FP_subtractor_13ccs_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_1 ( // @[FloatingPointDesigns.scala 1877:50]
    .clock(FP_subtractor_13ccs_1_clock),
    .reset(FP_subtractor_13ccs_1_reset),
    .io_in_a(FP_subtractor_13ccs_1_io_in_a),
    .io_in_b(FP_subtractor_13ccs_1_io_in_b),
    .io_out_s(FP_subtractor_13ccs_1_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_2 ( // @[FloatingPointDesigns.scala 1877:50]
    .clock(FP_subtractor_13ccs_2_clock),
    .reset(FP_subtractor_13ccs_2_reset),
    .io_in_a(FP_subtractor_13ccs_2_io_in_a),
    .io_in_b(FP_subtractor_13ccs_2_io_in_b),
    .io_out_s(FP_subtractor_13ccs_2_io_out_s)
  );
  FP_multiplier_10ccs multiplier4 ( // @[FloatingPointDesigns.scala 1945:29]
    .clock(multiplier4_clock),
    .reset(multiplier4_reset),
    .io_in_a(multiplier4_io_in_a),
    .io_in_b(multiplier4_io_in_b),
    .io_out_s(multiplier4_io_out_s)
  );
  assign io_out_s = {{1'd0}, multiplier4_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 1949:14]
  assign FP_multiplier_10ccs_clock = clock;
  assign FP_multiplier_10ccs_reset = reset;
  assign FP_multiplier_10ccs_io_in_a = {1'h0,result[30:0]}; // @[FloatingPointDesigns.scala 1903:48]
  assign FP_multiplier_10ccs_io_in_b = {1'h0,result[30:0]}; // @[FloatingPointDesigns.scala 1904:48]
  assign FP_multiplier_10ccs_1_clock = clock;
  assign FP_multiplier_10ccs_1_reset = reset;
  assign FP_multiplier_10ccs_1_io_in_a = FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 1916:34]
  assign FP_multiplier_10ccs_1_io_in_b = {1'h0,stage1_regs_0_1_8[30:0]}; // @[FloatingPointDesigns.scala 1917:46]
  assign FP_multiplier_10ccs_2_clock = clock;
  assign FP_multiplier_10ccs_2_reset = reset;
  assign FP_multiplier_10ccs_2_io_in_a = {1'h0,stage3_regs_0_0_11[30:0]}; // @[FloatingPointDesigns.scala 1934:46]
  assign FP_multiplier_10ccs_2_io_in_b = FP_subtractor_13ccs_io_out_s; // @[FloatingPointDesigns.scala 1935:34]
  assign FP_multiplier_10ccs_3_clock = clock;
  assign FP_multiplier_10ccs_3_reset = reset;
  assign FP_multiplier_10ccs_3_io_in_a = {1'h0,FP_multiplier_10ccs_2_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 1912:48]
  assign FP_multiplier_10ccs_3_io_in_b = {1'h0,FP_multiplier_10ccs_2_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 1913:48]
  assign FP_multiplier_10ccs_4_clock = clock;
  assign FP_multiplier_10ccs_4_reset = reset;
  assign FP_multiplier_10ccs_4_io_in_a = FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 1916:34]
  assign FP_multiplier_10ccs_4_io_in_b = {1'h0,stage1_regs_1_1_8[30:0]}; // @[FloatingPointDesigns.scala 1917:46]
  assign FP_multiplier_10ccs_5_clock = clock;
  assign FP_multiplier_10ccs_5_reset = reset;
  assign FP_multiplier_10ccs_5_io_in_a = {1'h0,stage3_regs_1_0_11[30:0]}; // @[FloatingPointDesigns.scala 1934:46]
  assign FP_multiplier_10ccs_5_io_in_b = FP_subtractor_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 1935:34]
  assign FP_multiplier_10ccs_6_clock = clock;
  assign FP_multiplier_10ccs_6_reset = reset;
  assign FP_multiplier_10ccs_6_io_in_a = {1'h0,FP_multiplier_10ccs_5_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 1912:48]
  assign FP_multiplier_10ccs_6_io_in_b = {1'h0,FP_multiplier_10ccs_5_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 1913:48]
  assign FP_multiplier_10ccs_7_clock = clock;
  assign FP_multiplier_10ccs_7_reset = reset;
  assign FP_multiplier_10ccs_7_io_in_a = FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 1916:34]
  assign FP_multiplier_10ccs_7_io_in_b = {1'h0,stage1_regs_2_1_8[30:0]}; // @[FloatingPointDesigns.scala 1917:46]
  assign FP_multiplier_10ccs_8_clock = clock;
  assign FP_multiplier_10ccs_8_reset = reset;
  assign FP_multiplier_10ccs_8_io_in_a = {1'h0,stage3_regs_2_0_11[30:0]}; // @[FloatingPointDesigns.scala 1934:46]
  assign FP_multiplier_10ccs_8_io_in_b = FP_subtractor_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 1935:34]
  assign FP_subtractor_13ccs_clock = clock;
  assign FP_subtractor_13ccs_reset = reset;
  assign FP_subtractor_13ccs_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1855:26 1856:16]
  assign FP_subtractor_13ccs_io_in_b = FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 1926:31]
  assign FP_subtractor_13ccs_1_clock = clock;
  assign FP_subtractor_13ccs_1_reset = reset;
  assign FP_subtractor_13ccs_1_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1855:26 1856:16]
  assign FP_subtractor_13ccs_1_io_in_b = FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 1926:31]
  assign FP_subtractor_13ccs_2_clock = clock;
  assign FP_subtractor_13ccs_2_reset = reset;
  assign FP_subtractor_13ccs_2_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1855:26 1856:16]
  assign FP_subtractor_13ccs_2_io_in_b = FP_multiplier_10ccs_7_io_out_s; // @[FloatingPointDesigns.scala 1926:31]
  assign multiplier4_clock = clock;
  assign multiplier4_reset = reset;
  assign multiplier4_io_in_a = {1'h0,FP_multiplier_10ccs_8_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 1947:37]
  assign multiplier4_io_in_b = {_restore_a_T_4,stage4_regs_2_1_8[22:0]}; // @[FloatingPointDesigns.scala 1944:113]
  always @(posedge clock) begin
    if (reset) begin // @[FloatingPointDesigns.scala 1869:22]
      x_n_0 <= 32'h0; // @[FloatingPointDesigns.scala 1869:22]
    end else begin
      x_n_0 <= result;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1869:22]
      x_n_1 <= 32'h0; // @[FloatingPointDesigns.scala 1869:22]
    end else begin
      x_n_1 <= stage1_regs_0_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1869:22]
      x_n_2 <= 32'h0; // @[FloatingPointDesigns.scala 1869:22]
    end else begin
      x_n_2 <= stage2_regs_0_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1869:22]
      x_n_4 <= 32'h0; // @[FloatingPointDesigns.scala 1869:22]
    end else begin
      x_n_4 <= _GEN_139;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1869:22]
      x_n_5 <= 32'h0; // @[FloatingPointDesigns.scala 1869:22]
    end else begin
      x_n_5 <= stage1_regs_1_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1869:22]
      x_n_6 <= 32'h0; // @[FloatingPointDesigns.scala 1869:22]
    end else begin
      x_n_6 <= stage2_regs_1_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1869:22]
      x_n_8 <= 32'h0; // @[FloatingPointDesigns.scala 1869:22]
    end else begin
      x_n_8 <= _GEN_215;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1869:22]
      x_n_9 <= 32'h0; // @[FloatingPointDesigns.scala 1869:22]
    end else begin
      x_n_9 <= stage1_regs_2_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1869:22]
      x_n_10 <= 32'h0; // @[FloatingPointDesigns.scala 1869:22]
    end else begin
      x_n_10 <= stage2_regs_2_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1870:22]
      a_2_0 <= 32'h0; // @[FloatingPointDesigns.scala 1870:22]
    end else begin
      a_2_0 <= _a_2_0_T_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1870:22]
      a_2_1 <= 32'h0; // @[FloatingPointDesigns.scala 1870:22]
    end else begin
      a_2_1 <= stage1_regs_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1870:22]
      a_2_2 <= 32'h0; // @[FloatingPointDesigns.scala 1870:22]
    end else begin
      a_2_2 <= stage2_regs_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1870:22]
      a_2_3 <= 32'h0; // @[FloatingPointDesigns.scala 1870:22]
    end else begin
      a_2_3 <= stage3_regs_0_1_11;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1870:22]
      a_2_4 <= 32'h0; // @[FloatingPointDesigns.scala 1870:22]
    end else begin
      a_2_4 <= stage4_regs_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1870:22]
      a_2_5 <= 32'h0; // @[FloatingPointDesigns.scala 1870:22]
    end else begin
      a_2_5 <= stage1_regs_1_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1870:22]
      a_2_6 <= 32'h0; // @[FloatingPointDesigns.scala 1870:22]
    end else begin
      a_2_6 <= stage2_regs_1_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1870:22]
      a_2_7 <= 32'h0; // @[FloatingPointDesigns.scala 1870:22]
    end else begin
      a_2_7 <= stage3_regs_1_1_11;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1870:22]
      a_2_8 <= 32'h0; // @[FloatingPointDesigns.scala 1870:22]
    end else begin
      a_2_8 <= stage4_regs_1_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1870:22]
      a_2_9 <= 32'h0; // @[FloatingPointDesigns.scala 1870:22]
    end else begin
      a_2_9 <= stage1_regs_2_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1870:22]
      a_2_10 <= 32'h0; // @[FloatingPointDesigns.scala 1870:22]
    end else begin
      a_2_10 <= stage2_regs_2_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1870:22]
      a_2_11 <= 32'h0; // @[FloatingPointDesigns.scala 1870:22]
    end else begin
      a_2_11 <= stage3_regs_2_1_11;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_0_0 <= x_n_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_0_1 <= stage1_regs_0_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_0_2 <= stage1_regs_0_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_0_3 <= stage1_regs_0_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_0_4 <= stage1_regs_0_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_0_5 <= stage1_regs_0_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_0_6 <= stage1_regs_0_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_0_7 <= stage1_regs_0_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_0_8 <= stage1_regs_0_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_1_0 <= a_2_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_1_1 <= stage1_regs_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_1_2 <= stage1_regs_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_1_3 <= stage1_regs_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_1_4 <= stage1_regs_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_1_5 <= stage1_regs_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_1_6 <= stage1_regs_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_1_7 <= stage1_regs_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_0_1_8 <= stage1_regs_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_0_0 <= x_n_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_0_1 <= stage1_regs_1_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_0_2 <= stage1_regs_1_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_0_3 <= stage1_regs_1_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_0_4 <= stage1_regs_1_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_0_5 <= stage1_regs_1_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_0_6 <= stage1_regs_1_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_0_7 <= stage1_regs_1_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_0_8 <= stage1_regs_1_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_1_0 <= a_2_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_1_1 <= stage1_regs_1_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_1_2 <= stage1_regs_1_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_1_3 <= stage1_regs_1_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_1_4 <= stage1_regs_1_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_1_5 <= stage1_regs_1_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_1_6 <= stage1_regs_1_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_1_7 <= stage1_regs_1_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_1_1_8 <= stage1_regs_1_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_0_0 <= x_n_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_0_1 <= stage1_regs_2_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_0_2 <= stage1_regs_2_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_0_3 <= stage1_regs_2_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_0_4 <= stage1_regs_2_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_0_5 <= stage1_regs_2_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_0_6 <= stage1_regs_2_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_0_7 <= stage1_regs_2_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_0_8 <= stage1_regs_2_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_1_0 <= a_2_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_1_1 <= stage1_regs_2_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_1_2 <= stage1_regs_2_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_1_3 <= stage1_regs_2_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_1_4 <= stage1_regs_2_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_1_5 <= stage1_regs_2_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_1_6 <= stage1_regs_2_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_1_7 <= stage1_regs_2_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:30]
      stage1_regs_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1871:30]
    end else begin
      stage1_regs_2_1_8 <= stage1_regs_2_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_0_0 <= x_n_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_0_1 <= stage2_regs_0_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_0_2 <= stage2_regs_0_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_0_3 <= stage2_regs_0_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_0_4 <= stage2_regs_0_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_0_5 <= stage2_regs_0_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_0_6 <= stage2_regs_0_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_0_7 <= stage2_regs_0_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_0_8 <= stage2_regs_0_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_1_0 <= a_2_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_1_1 <= stage2_regs_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_1_2 <= stage2_regs_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_1_3 <= stage2_regs_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_1_4 <= stage2_regs_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_1_5 <= stage2_regs_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_1_6 <= stage2_regs_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_1_7 <= stage2_regs_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_0_1_8 <= stage2_regs_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_0_0 <= x_n_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_0_1 <= stage2_regs_1_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_0_2 <= stage2_regs_1_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_0_3 <= stage2_regs_1_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_0_4 <= stage2_regs_1_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_0_5 <= stage2_regs_1_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_0_6 <= stage2_regs_1_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_0_7 <= stage2_regs_1_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_0_8 <= stage2_regs_1_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_1_0 <= a_2_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_1_1 <= stage2_regs_1_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_1_2 <= stage2_regs_1_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_1_3 <= stage2_regs_1_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_1_4 <= stage2_regs_1_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_1_5 <= stage2_regs_1_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_1_6 <= stage2_regs_1_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_1_7 <= stage2_regs_1_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_1_1_8 <= stage2_regs_1_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_0_0 <= x_n_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_0_1 <= stage2_regs_2_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_0_2 <= stage2_regs_2_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_0_3 <= stage2_regs_2_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_0_4 <= stage2_regs_2_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_0_5 <= stage2_regs_2_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_0_6 <= stage2_regs_2_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_0_7 <= stage2_regs_2_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_0_8 <= stage2_regs_2_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_1_0 <= a_2_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_1_1 <= stage2_regs_2_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_1_2 <= stage2_regs_2_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_1_3 <= stage2_regs_2_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_1_4 <= stage2_regs_2_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_1_5 <= stage2_regs_2_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_1_6 <= stage2_regs_2_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_1_7 <= stage2_regs_2_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:30]
      stage2_regs_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1872:30]
    end else begin
      stage2_regs_2_1_8 <= stage2_regs_2_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_0_0 <= x_n_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_0_1 <= stage3_regs_0_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_0_2 <= stage3_regs_0_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_0_3 <= stage3_regs_0_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_0_4 <= stage3_regs_0_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_0_5 <= stage3_regs_0_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_0_6 <= stage3_regs_0_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_0_7 <= stage3_regs_0_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_0_8 <= stage3_regs_0_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_0_9 <= stage3_regs_0_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_0_10 <= stage3_regs_0_0_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_0_11 <= stage3_regs_0_0_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_1_0 <= a_2_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_1_1 <= stage3_regs_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_1_2 <= stage3_regs_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_1_3 <= stage3_regs_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_1_4 <= stage3_regs_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_1_5 <= stage3_regs_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_1_6 <= stage3_regs_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_1_7 <= stage3_regs_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_1_8 <= stage3_regs_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_1_9 <= stage3_regs_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_1_10 <= stage3_regs_0_1_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_0_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_0_1_11 <= stage3_regs_0_1_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_0_0 <= x_n_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_0_1 <= stage3_regs_1_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_0_2 <= stage3_regs_1_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_0_3 <= stage3_regs_1_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_0_4 <= stage3_regs_1_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_0_5 <= stage3_regs_1_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_0_6 <= stage3_regs_1_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_0_7 <= stage3_regs_1_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_0_8 <= stage3_regs_1_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_0_9 <= stage3_regs_1_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_0_10 <= stage3_regs_1_0_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_0_11 <= stage3_regs_1_0_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_1_0 <= a_2_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_1_1 <= stage3_regs_1_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_1_2 <= stage3_regs_1_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_1_3 <= stage3_regs_1_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_1_4 <= stage3_regs_1_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_1_5 <= stage3_regs_1_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_1_6 <= stage3_regs_1_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_1_7 <= stage3_regs_1_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_1_8 <= stage3_regs_1_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_1_9 <= stage3_regs_1_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_1_10 <= stage3_regs_1_1_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_1_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_1_1_11 <= stage3_regs_1_1_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_0_0 <= x_n_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_0_1 <= stage3_regs_2_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_0_2 <= stage3_regs_2_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_0_3 <= stage3_regs_2_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_0_4 <= stage3_regs_2_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_0_5 <= stage3_regs_2_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_0_6 <= stage3_regs_2_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_0_7 <= stage3_regs_2_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_0_8 <= stage3_regs_2_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_0_9 <= stage3_regs_2_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_0_10 <= stage3_regs_2_0_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_0_11 <= stage3_regs_2_0_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_1_0 <= a_2_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_1_1 <= stage3_regs_2_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_1_2 <= stage3_regs_2_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_1_3 <= stage3_regs_2_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_1_4 <= stage3_regs_2_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_1_5 <= stage3_regs_2_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_1_6 <= stage3_regs_2_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_1_7 <= stage3_regs_2_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_1_8 <= stage3_regs_2_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_1_9 <= stage3_regs_2_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_1_10 <= stage3_regs_2_1_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage3_regs_2_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage3_regs_2_1_11 <= stage3_regs_2_1_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_0_1_0 <= a_2_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_0_1_1 <= stage4_regs_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_0_1_2 <= stage4_regs_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_0_1_3 <= stage4_regs_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_0_1_4 <= stage4_regs_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_0_1_5 <= stage4_regs_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_0_1_6 <= stage4_regs_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_0_1_7 <= stage4_regs_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_0_1_8 <= stage4_regs_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_1_1_0 <= a_2_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_1_1_1 <= stage4_regs_1_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_1_1_2 <= stage4_regs_1_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_1_1_3 <= stage4_regs_1_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_1_1_4 <= stage4_regs_1_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_1_1_5 <= stage4_regs_1_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_1_1_6 <= stage4_regs_1_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_1_1_7 <= stage4_regs_1_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_1_1_8 <= stage4_regs_1_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_2_1_0 <= a_2_11;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_2_1_1 <= stage4_regs_2_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_2_1_2 <= stage4_regs_2_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_2_1_3 <= stage4_regs_2_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_2_1_4 <= stage4_regs_2_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_2_1_5 <= stage4_regs_2_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_2_1_6 <= stage4_regs_2_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_2_1_7 <= stage4_regs_2_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage4_regs_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage4_regs_2_1_8 <= stage4_regs_2_1_7;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  x_n_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  x_n_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  x_n_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  x_n_4 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  x_n_5 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  x_n_6 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  x_n_8 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  x_n_9 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  x_n_10 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  a_2_0 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  a_2_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  a_2_2 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  a_2_3 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  a_2_4 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  a_2_5 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  a_2_6 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  a_2_7 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  a_2_8 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  a_2_9 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  a_2_10 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  a_2_11 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  stage1_regs_0_0_0 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  stage1_regs_0_0_1 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  stage1_regs_0_0_2 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  stage1_regs_0_0_3 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  stage1_regs_0_0_4 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  stage1_regs_0_0_5 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  stage1_regs_0_0_6 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  stage1_regs_0_0_7 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  stage1_regs_0_0_8 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  stage1_regs_0_1_0 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  stage1_regs_0_1_1 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  stage1_regs_0_1_2 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  stage1_regs_0_1_3 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  stage1_regs_0_1_4 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  stage1_regs_0_1_5 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  stage1_regs_0_1_6 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  stage1_regs_0_1_7 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  stage1_regs_0_1_8 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  stage1_regs_1_0_0 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  stage1_regs_1_0_1 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  stage1_regs_1_0_2 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  stage1_regs_1_0_3 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  stage1_regs_1_0_4 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  stage1_regs_1_0_5 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  stage1_regs_1_0_6 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  stage1_regs_1_0_7 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  stage1_regs_1_0_8 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  stage1_regs_1_1_0 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  stage1_regs_1_1_1 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  stage1_regs_1_1_2 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  stage1_regs_1_1_3 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  stage1_regs_1_1_4 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  stage1_regs_1_1_5 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  stage1_regs_1_1_6 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  stage1_regs_1_1_7 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  stage1_regs_1_1_8 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  stage1_regs_2_0_0 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  stage1_regs_2_0_1 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  stage1_regs_2_0_2 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  stage1_regs_2_0_3 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  stage1_regs_2_0_4 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  stage1_regs_2_0_5 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  stage1_regs_2_0_6 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  stage1_regs_2_0_7 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  stage1_regs_2_0_8 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  stage1_regs_2_1_0 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  stage1_regs_2_1_1 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  stage1_regs_2_1_2 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  stage1_regs_2_1_3 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  stage1_regs_2_1_4 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  stage1_regs_2_1_5 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  stage1_regs_2_1_6 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  stage1_regs_2_1_7 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  stage1_regs_2_1_8 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  stage2_regs_0_0_0 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  stage2_regs_0_0_1 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  stage2_regs_0_0_2 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  stage2_regs_0_0_3 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  stage2_regs_0_0_4 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  stage2_regs_0_0_5 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  stage2_regs_0_0_6 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  stage2_regs_0_0_7 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  stage2_regs_0_0_8 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  stage2_regs_0_1_0 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  stage2_regs_0_1_1 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  stage2_regs_0_1_2 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  stage2_regs_0_1_3 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  stage2_regs_0_1_4 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  stage2_regs_0_1_5 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  stage2_regs_0_1_6 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  stage2_regs_0_1_7 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  stage2_regs_0_1_8 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  stage2_regs_1_0_0 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  stage2_regs_1_0_1 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  stage2_regs_1_0_2 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  stage2_regs_1_0_3 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  stage2_regs_1_0_4 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  stage2_regs_1_0_5 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  stage2_regs_1_0_6 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  stage2_regs_1_0_7 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  stage2_regs_1_0_8 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  stage2_regs_1_1_0 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  stage2_regs_1_1_1 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  stage2_regs_1_1_2 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  stage2_regs_1_1_3 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  stage2_regs_1_1_4 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  stage2_regs_1_1_5 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  stage2_regs_1_1_6 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  stage2_regs_1_1_7 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  stage2_regs_1_1_8 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  stage2_regs_2_0_0 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  stage2_regs_2_0_1 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  stage2_regs_2_0_2 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  stage2_regs_2_0_3 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  stage2_regs_2_0_4 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  stage2_regs_2_0_5 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  stage2_regs_2_0_6 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  stage2_regs_2_0_7 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  stage2_regs_2_0_8 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  stage2_regs_2_1_0 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  stage2_regs_2_1_1 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  stage2_regs_2_1_2 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  stage2_regs_2_1_3 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  stage2_regs_2_1_4 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  stage2_regs_2_1_5 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  stage2_regs_2_1_6 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  stage2_regs_2_1_7 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  stage2_regs_2_1_8 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  stage3_regs_0_0_0 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  stage3_regs_0_0_1 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  stage3_regs_0_0_2 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  stage3_regs_0_0_3 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  stage3_regs_0_0_4 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  stage3_regs_0_0_5 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  stage3_regs_0_0_6 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  stage3_regs_0_0_7 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  stage3_regs_0_0_8 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  stage3_regs_0_0_9 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  stage3_regs_0_0_10 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  stage3_regs_0_0_11 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  stage3_regs_0_1_0 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  stage3_regs_0_1_1 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  stage3_regs_0_1_2 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  stage3_regs_0_1_3 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  stage3_regs_0_1_4 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  stage3_regs_0_1_5 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  stage3_regs_0_1_6 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  stage3_regs_0_1_7 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  stage3_regs_0_1_8 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  stage3_regs_0_1_9 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  stage3_regs_0_1_10 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  stage3_regs_0_1_11 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  stage3_regs_1_0_0 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  stage3_regs_1_0_1 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  stage3_regs_1_0_2 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  stage3_regs_1_0_3 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  stage3_regs_1_0_4 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  stage3_regs_1_0_5 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  stage3_regs_1_0_6 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  stage3_regs_1_0_7 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  stage3_regs_1_0_8 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  stage3_regs_1_0_9 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  stage3_regs_1_0_10 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  stage3_regs_1_0_11 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  stage3_regs_1_1_0 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  stage3_regs_1_1_1 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  stage3_regs_1_1_2 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  stage3_regs_1_1_3 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  stage3_regs_1_1_4 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  stage3_regs_1_1_5 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  stage3_regs_1_1_6 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  stage3_regs_1_1_7 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  stage3_regs_1_1_8 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  stage3_regs_1_1_9 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  stage3_regs_1_1_10 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  stage3_regs_1_1_11 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  stage3_regs_2_0_0 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  stage3_regs_2_0_1 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  stage3_regs_2_0_2 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  stage3_regs_2_0_3 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  stage3_regs_2_0_4 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  stage3_regs_2_0_5 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  stage3_regs_2_0_6 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  stage3_regs_2_0_7 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  stage3_regs_2_0_8 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  stage3_regs_2_0_9 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  stage3_regs_2_0_10 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  stage3_regs_2_0_11 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  stage3_regs_2_1_0 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  stage3_regs_2_1_1 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  stage3_regs_2_1_2 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  stage3_regs_2_1_3 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  stage3_regs_2_1_4 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  stage3_regs_2_1_5 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  stage3_regs_2_1_6 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  stage3_regs_2_1_7 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  stage3_regs_2_1_8 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  stage3_regs_2_1_9 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  stage3_regs_2_1_10 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  stage3_regs_2_1_11 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  stage4_regs_0_1_0 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  stage4_regs_0_1_1 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  stage4_regs_0_1_2 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  stage4_regs_0_1_3 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  stage4_regs_0_1_4 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  stage4_regs_0_1_5 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  stage4_regs_0_1_6 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  stage4_regs_0_1_7 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  stage4_regs_0_1_8 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  stage4_regs_1_1_0 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  stage4_regs_1_1_1 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  stage4_regs_1_1_2 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  stage4_regs_1_1_3 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  stage4_regs_1_1_4 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  stage4_regs_1_1_5 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  stage4_regs_1_1_6 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  stage4_regs_1_1_7 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  stage4_regs_1_1_8 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  stage4_regs_2_1_0 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  stage4_regs_2_1_1 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  stage4_regs_2_1_2 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  stage4_regs_2_1_3 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  stage4_regs_2_1_4 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  stage4_regs_2_1_5 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  stage4_regs_2_1_6 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  stage4_regs_2_1_7 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  stage4_regs_2_1_8 = _RAND_227[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module hqr5(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
  wire  FP_adder_13ccs_clock; // @[FloatingPointDesigns.scala 2510:23]
  wire  FP_adder_13ccs_reset; // @[FloatingPointDesigns.scala 2510:23]
  wire [31:0] FP_adder_13ccs_io_in_a; // @[FloatingPointDesigns.scala 2510:23]
  wire [31:0] FP_adder_13ccs_io_in_b; // @[FloatingPointDesigns.scala 2510:23]
  wire [31:0] FP_adder_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2510:23]
  wire  FP_subtractor_13ccs_clock; // @[FloatingPointDesigns.scala 2511:28]
  wire  FP_subtractor_13ccs_reset; // @[FloatingPointDesigns.scala 2511:28]
  wire [31:0] FP_subtractor_13ccs_io_in_a; // @[FloatingPointDesigns.scala 2511:28]
  wire [31:0] FP_subtractor_13ccs_io_in_b; // @[FloatingPointDesigns.scala 2511:28]
  wire [31:0] FP_subtractor_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2511:28]
  FP_adder_13ccs FP_adder_13ccs ( // @[FloatingPointDesigns.scala 2510:23]
    .clock(FP_adder_13ccs_clock),
    .reset(FP_adder_13ccs_reset),
    .io_in_a(FP_adder_13ccs_io_in_a),
    .io_in_b(FP_adder_13ccs_io_in_b),
    .io_out_s(FP_adder_13ccs_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs ( // @[FloatingPointDesigns.scala 2511:28]
    .clock(FP_subtractor_13ccs_clock),
    .reset(FP_subtractor_13ccs_reset),
    .io_in_a(FP_subtractor_13ccs_io_in_a),
    .io_in_b(FP_subtractor_13ccs_io_in_b),
    .io_out_s(FP_subtractor_13ccs_io_out_s)
  );
  assign io_out_s = io_in_a[31] ? FP_subtractor_13ccs_io_out_s : FP_adder_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2519:24 2520:14 2522:14]
  assign FP_adder_13ccs_clock = clock;
  assign FP_adder_13ccs_reset = reset;
  assign FP_adder_13ccs_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2513:16]
  assign FP_adder_13ccs_io_in_b = io_in_b; // @[FloatingPointDesigns.scala 2514:16]
  assign FP_subtractor_13ccs_clock = clock;
  assign FP_subtractor_13ccs_reset = reset;
  assign FP_subtractor_13ccs_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2516:21]
  assign FP_subtractor_13ccs_io_in_b = io_in_b; // @[FloatingPointDesigns.scala 2517:21]
endmodule
module FP_reciprocal_newfpu(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
`endif // RANDOMIZE_REG_INIT
  wire  FP_multiplier_10ccs_clock; // @[FloatingPointDesigns.scala 2005:65]
  wire  FP_multiplier_10ccs_reset; // @[FloatingPointDesigns.scala 2005:65]
  wire [31:0] FP_multiplier_10ccs_io_in_a; // @[FloatingPointDesigns.scala 2005:65]
  wire [31:0] FP_multiplier_10ccs_io_in_b; // @[FloatingPointDesigns.scala 2005:65]
  wire [31:0] FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2005:65]
  wire  FP_multiplier_10ccs_1_clock; // @[FloatingPointDesigns.scala 2005:65]
  wire  FP_multiplier_10ccs_1_reset; // @[FloatingPointDesigns.scala 2005:65]
  wire [31:0] FP_multiplier_10ccs_1_io_in_a; // @[FloatingPointDesigns.scala 2005:65]
  wire [31:0] FP_multiplier_10ccs_1_io_in_b; // @[FloatingPointDesigns.scala 2005:65]
  wire [31:0] FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2005:65]
  wire  FP_multiplier_10ccs_2_clock; // @[FloatingPointDesigns.scala 2005:65]
  wire  FP_multiplier_10ccs_2_reset; // @[FloatingPointDesigns.scala 2005:65]
  wire [31:0] FP_multiplier_10ccs_2_io_in_a; // @[FloatingPointDesigns.scala 2005:65]
  wire [31:0] FP_multiplier_10ccs_2_io_in_b; // @[FloatingPointDesigns.scala 2005:65]
  wire [31:0] FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2005:65]
  wire  FP_subtractor_13ccs_clock; // @[FloatingPointDesigns.scala 2006:50]
  wire  FP_subtractor_13ccs_reset; // @[FloatingPointDesigns.scala 2006:50]
  wire [31:0] FP_subtractor_13ccs_io_in_a; // @[FloatingPointDesigns.scala 2006:50]
  wire [31:0] FP_subtractor_13ccs_io_in_b; // @[FloatingPointDesigns.scala 2006:50]
  wire [31:0] FP_subtractor_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2006:50]
  wire  multiplier4_clock; // @[FloatingPointDesigns.scala 2085:29]
  wire  multiplier4_reset; // @[FloatingPointDesigns.scala 2085:29]
  wire [31:0] multiplier4_io_in_a; // @[FloatingPointDesigns.scala 2085:29]
  wire [31:0] multiplier4_io_in_b; // @[FloatingPointDesigns.scala 2085:29]
  wire [31:0] multiplier4_io_out_s; // @[FloatingPointDesigns.scala 2085:29]
  wire  FP_multiplier_10ccs_3_clock; // @[FloatingPointDesigns.scala 2097:69]
  wire  FP_multiplier_10ccs_3_reset; // @[FloatingPointDesigns.scala 2097:69]
  wire [31:0] FP_multiplier_10ccs_3_io_in_a; // @[FloatingPointDesigns.scala 2097:69]
  wire [31:0] FP_multiplier_10ccs_3_io_in_b; // @[FloatingPointDesigns.scala 2097:69]
  wire [31:0] FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2097:69]
  wire  FP_multiplier_10ccs_4_clock; // @[FloatingPointDesigns.scala 2097:69]
  wire  FP_multiplier_10ccs_4_reset; // @[FloatingPointDesigns.scala 2097:69]
  wire [31:0] FP_multiplier_10ccs_4_io_in_a; // @[FloatingPointDesigns.scala 2097:69]
  wire [31:0] FP_multiplier_10ccs_4_io_in_b; // @[FloatingPointDesigns.scala 2097:69]
  wire [31:0] FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2097:69]
  wire  FP_multiplier_10ccs_5_clock; // @[FloatingPointDesigns.scala 2097:69]
  wire  FP_multiplier_10ccs_5_reset; // @[FloatingPointDesigns.scala 2097:69]
  wire [31:0] FP_multiplier_10ccs_5_io_in_a; // @[FloatingPointDesigns.scala 2097:69]
  wire [31:0] FP_multiplier_10ccs_5_io_in_b; // @[FloatingPointDesigns.scala 2097:69]
  wire [31:0] FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2097:69]
  wire  FP_multiplier_10ccs_6_clock; // @[FloatingPointDesigns.scala 2097:69]
  wire  FP_multiplier_10ccs_6_reset; // @[FloatingPointDesigns.scala 2097:69]
  wire [31:0] FP_multiplier_10ccs_6_io_in_a; // @[FloatingPointDesigns.scala 2097:69]
  wire [31:0] FP_multiplier_10ccs_6_io_in_b; // @[FloatingPointDesigns.scala 2097:69]
  wire [31:0] FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2097:69]
  wire  FP_subtractor_13ccs_1_clock; // @[FloatingPointDesigns.scala 2098:54]
  wire  FP_subtractor_13ccs_1_reset; // @[FloatingPointDesigns.scala 2098:54]
  wire [31:0] FP_subtractor_13ccs_1_io_in_a; // @[FloatingPointDesigns.scala 2098:54]
  wire [31:0] FP_subtractor_13ccs_1_io_in_b; // @[FloatingPointDesigns.scala 2098:54]
  wire [31:0] FP_subtractor_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2098:54]
  wire  FP_subtractor_13ccs_2_clock; // @[FloatingPointDesigns.scala 2098:54]
  wire  FP_subtractor_13ccs_2_reset; // @[FloatingPointDesigns.scala 2098:54]
  wire [31:0] FP_subtractor_13ccs_2_io_in_a; // @[FloatingPointDesigns.scala 2098:54]
  wire [31:0] FP_subtractor_13ccs_2_io_in_b; // @[FloatingPointDesigns.scala 2098:54]
  wire [31:0] FP_subtractor_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2098:54]
  wire [30:0] _number_T_1 = {{1'd0}, io_in_a[30:1]}; // @[FloatingPointDesigns.scala 1990:36]
  wire [30:0] _GEN_0 = io_in_a[30:0] > 31'h7ef477d4 ? 31'h3f7a3bea : _number_T_1; // @[FloatingPointDesigns.scala 1987:46 1988:14 1990:14]
  wire [31:0] number = {{1'd0}, _GEN_0}; // @[FloatingPointDesigns.scala 1982:22]
  wire [31:0] result = 32'h5f3759df - number; // @[FloatingPointDesigns.scala 1997:25]
  reg [31:0] x_n_0; // @[FloatingPointDesigns.scala 1999:22]
  reg [31:0] x_n_1; // @[FloatingPointDesigns.scala 1999:22]
  reg [31:0] x_n_2; // @[FloatingPointDesigns.scala 1999:22]
  reg [31:0] a_2_0; // @[FloatingPointDesigns.scala 2000:22]
  reg [31:0] a_2_1; // @[FloatingPointDesigns.scala 2000:22]
  reg [31:0] a_2_2; // @[FloatingPointDesigns.scala 2000:22]
  reg [31:0] a_2_3; // @[FloatingPointDesigns.scala 2000:22]
  reg [31:0] stage1_regs_0_0_0; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage1_regs_0_0_1; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage1_regs_0_0_2; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage1_regs_0_0_3; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage1_regs_0_0_4; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage1_regs_0_0_5; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage1_regs_0_0_6; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage1_regs_0_0_7; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage1_regs_0_0_8; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage1_regs_0_1_0; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage1_regs_0_1_1; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage1_regs_0_1_2; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage1_regs_0_1_3; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage1_regs_0_1_4; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage1_regs_0_1_5; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage1_regs_0_1_6; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage1_regs_0_1_7; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage1_regs_0_1_8; // @[FloatingPointDesigns.scala 2001:30]
  reg [31:0] stage2_regs_0_0_0; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage2_regs_0_0_1; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage2_regs_0_0_2; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage2_regs_0_0_3; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage2_regs_0_0_4; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage2_regs_0_0_5; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage2_regs_0_0_6; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage2_regs_0_0_7; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage2_regs_0_0_8; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage2_regs_0_1_0; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage2_regs_0_1_1; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage2_regs_0_1_2; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage2_regs_0_1_3; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage2_regs_0_1_4; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage2_regs_0_1_5; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage2_regs_0_1_6; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage2_regs_0_1_7; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage2_regs_0_1_8; // @[FloatingPointDesigns.scala 2002:30]
  reg [31:0] stage3_regs_0_0_0; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_0_1; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_0_2; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_0_3; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_0_4; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_0_5; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_0_6; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_0_7; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_0_8; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_0_9; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_0_10; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_0_11; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_1_0; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_1_1; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_1_2; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_1_3; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_1_4; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_1_5; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_1_6; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_1_7; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_1_8; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_1_9; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_1_10; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage3_regs_0_1_11; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage4_regs_0_1_0; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage4_regs_0_1_1; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage4_regs_0_1_2; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage4_regs_0_1_3; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage4_regs_0_1_4; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage4_regs_0_1_5; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage4_regs_0_1_6; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage4_regs_0_1_7; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage4_regs_0_1_8; // @[FloatingPointDesigns.scala 2004:30]
  wire [7:0] _a_2_0_T_3 = io_in_a[30:23] - 8'h1; // @[FloatingPointDesigns.scala 2030:75]
  wire [31:0] _a_2_0_T_6 = {io_in_a[31],_a_2_0_T_3,io_in_a[22:0]}; // @[FloatingPointDesigns.scala 2030:82]
  reg [31:0] a_2_isr_to_r; // @[FloatingPointDesigns.scala 2075:31]
  reg [31:0] transition_regs_0; // @[FloatingPointDesigns.scala 2076:34]
  reg [31:0] transition_regs_1; // @[FloatingPointDesigns.scala 2076:34]
  reg [31:0] transition_regs_2; // @[FloatingPointDesigns.scala 2076:34]
  reg [31:0] transition_regs_3; // @[FloatingPointDesigns.scala 2076:34]
  reg [31:0] transition_regs_4; // @[FloatingPointDesigns.scala 2076:34]
  reg [31:0] transition_regs_5; // @[FloatingPointDesigns.scala 2076:34]
  reg [31:0] transition_regs_6; // @[FloatingPointDesigns.scala 2076:34]
  reg [31:0] transition_regs_7; // @[FloatingPointDesigns.scala 2076:34]
  reg [31:0] transition_regs_8; // @[FloatingPointDesigns.scala 2076:34]
  wire [7:0] _a_2_isr_to_r_T_3 = stage4_regs_0_1_8[30:23] + 8'h1; // @[FloatingPointDesigns.scala 2078:115]
  wire [31:0] _a_2_isr_to_r_T_6 = {stage4_regs_0_1_8[31],_a_2_isr_to_r_T_3,stage4_regs_0_1_8[22:0]}; // @[FloatingPointDesigns.scala 2078:122]
  reg [31:0] x_n_r_0; // @[FloatingPointDesigns.scala 2092:24]
  reg [31:0] x_n_r_1; // @[FloatingPointDesigns.scala 2092:24]
  reg [31:0] x_n_r_3; // @[FloatingPointDesigns.scala 2092:24]
  reg [31:0] x_n_r_4; // @[FloatingPointDesigns.scala 2092:24]
  reg [31:0] a_2_r_0; // @[FloatingPointDesigns.scala 2093:24]
  reg [31:0] a_2_r_1; // @[FloatingPointDesigns.scala 2093:24]
  reg [31:0] a_2_r_2; // @[FloatingPointDesigns.scala 2093:24]
  reg [31:0] a_2_r_3; // @[FloatingPointDesigns.scala 2093:24]
  reg [31:0] a_2_r_4; // @[FloatingPointDesigns.scala 2093:24]
  reg [31:0] a_2_r_5; // @[FloatingPointDesigns.scala 2093:24]
  reg [31:0] stage1_regs_r_0_0_0; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_0_0_1; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_0_0_2; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_0_0_3; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_0_0_4; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_0_0_5; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_0_0_6; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_0_0_7; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_0_0_8; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_0_1_0; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_0_1_1; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_0_1_2; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_0_1_3; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_0_1_4; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_0_1_5; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_0_1_6; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_0_1_7; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_0_1_8; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_0_0; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_0_1; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_0_2; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_0_3; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_0_4; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_0_5; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_0_6; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_0_7; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_0_8; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_1_0; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_1_1; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_1_2; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_1_3; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_1_4; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_1_5; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_1_6; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_1_7; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage1_regs_r_1_1_8; // @[FloatingPointDesigns.scala 2094:32]
  reg [31:0] stage2_regs_r_0_0_0; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_0_1; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_0_2; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_0_3; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_0_4; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_0_5; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_0_6; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_0_7; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_0_8; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_0_9; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_0_10; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_0_11; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_1_0; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_1_1; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_1_2; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_1_3; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_1_4; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_1_5; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_1_6; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_1_7; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_1_8; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_1_9; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_1_10; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_0_1_11; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_0_0; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_0_1; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_0_2; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_0_3; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_0_4; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_0_5; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_0_6; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_0_7; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_0_8; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_0_9; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_0_10; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_0_11; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_1_0; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_1_1; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_1_2; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_1_3; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_1_4; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_1_5; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_1_6; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_1_7; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_1_8; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_1_9; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_1_10; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage2_regs_r_1_1_11; // @[FloatingPointDesigns.scala 2095:32]
  reg [31:0] stage3_regs_r_0_1_0; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage3_regs_r_0_1_1; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage3_regs_r_0_1_2; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage3_regs_r_0_1_3; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage3_regs_r_0_1_4; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage3_regs_r_0_1_5; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage3_regs_r_0_1_6; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage3_regs_r_0_1_7; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage3_regs_r_0_1_8; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage3_regs_r_1_1_0; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage3_regs_r_1_1_1; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage3_regs_r_1_1_2; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage3_regs_r_1_1_3; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage3_regs_r_1_1_4; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage3_regs_r_1_1_5; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage3_regs_r_1_1_6; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage3_regs_r_1_1_7; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage3_regs_r_1_1_8; // @[FloatingPointDesigns.scala 2096:32]
  wire [31:0] _GEN_133 = multiplier4_io_out_s; // @[FloatingPointDesigns.scala 2092:24 2117:28 2118:28]
  wire [31:0] _GEN_189 = FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2092:24 2126:28 2127:28]
  FP_multiplier_10ccs FP_multiplier_10ccs ( // @[FloatingPointDesigns.scala 2005:65]
    .clock(FP_multiplier_10ccs_clock),
    .reset(FP_multiplier_10ccs_reset),
    .io_in_a(FP_multiplier_10ccs_io_in_a),
    .io_in_b(FP_multiplier_10ccs_io_in_b),
    .io_out_s(FP_multiplier_10ccs_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_1 ( // @[FloatingPointDesigns.scala 2005:65]
    .clock(FP_multiplier_10ccs_1_clock),
    .reset(FP_multiplier_10ccs_1_reset),
    .io_in_a(FP_multiplier_10ccs_1_io_in_a),
    .io_in_b(FP_multiplier_10ccs_1_io_in_b),
    .io_out_s(FP_multiplier_10ccs_1_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_2 ( // @[FloatingPointDesigns.scala 2005:65]
    .clock(FP_multiplier_10ccs_2_clock),
    .reset(FP_multiplier_10ccs_2_reset),
    .io_in_a(FP_multiplier_10ccs_2_io_in_a),
    .io_in_b(FP_multiplier_10ccs_2_io_in_b),
    .io_out_s(FP_multiplier_10ccs_2_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs ( // @[FloatingPointDesigns.scala 2006:50]
    .clock(FP_subtractor_13ccs_clock),
    .reset(FP_subtractor_13ccs_reset),
    .io_in_a(FP_subtractor_13ccs_io_in_a),
    .io_in_b(FP_subtractor_13ccs_io_in_b),
    .io_out_s(FP_subtractor_13ccs_io_out_s)
  );
  FP_multiplier_10ccs multiplier4 ( // @[FloatingPointDesigns.scala 2085:29]
    .clock(multiplier4_clock),
    .reset(multiplier4_reset),
    .io_in_a(multiplier4_io_in_a),
    .io_in_b(multiplier4_io_in_b),
    .io_out_s(multiplier4_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_3 ( // @[FloatingPointDesigns.scala 2097:69]
    .clock(FP_multiplier_10ccs_3_clock),
    .reset(FP_multiplier_10ccs_3_reset),
    .io_in_a(FP_multiplier_10ccs_3_io_in_a),
    .io_in_b(FP_multiplier_10ccs_3_io_in_b),
    .io_out_s(FP_multiplier_10ccs_3_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_4 ( // @[FloatingPointDesigns.scala 2097:69]
    .clock(FP_multiplier_10ccs_4_clock),
    .reset(FP_multiplier_10ccs_4_reset),
    .io_in_a(FP_multiplier_10ccs_4_io_in_a),
    .io_in_b(FP_multiplier_10ccs_4_io_in_b),
    .io_out_s(FP_multiplier_10ccs_4_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_5 ( // @[FloatingPointDesigns.scala 2097:69]
    .clock(FP_multiplier_10ccs_5_clock),
    .reset(FP_multiplier_10ccs_5_reset),
    .io_in_a(FP_multiplier_10ccs_5_io_in_a),
    .io_in_b(FP_multiplier_10ccs_5_io_in_b),
    .io_out_s(FP_multiplier_10ccs_5_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_6 ( // @[FloatingPointDesigns.scala 2097:69]
    .clock(FP_multiplier_10ccs_6_clock),
    .reset(FP_multiplier_10ccs_6_reset),
    .io_in_a(FP_multiplier_10ccs_6_io_in_a),
    .io_in_b(FP_multiplier_10ccs_6_io_in_b),
    .io_out_s(FP_multiplier_10ccs_6_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_1 ( // @[FloatingPointDesigns.scala 2098:54]
    .clock(FP_subtractor_13ccs_1_clock),
    .reset(FP_subtractor_13ccs_1_reset),
    .io_in_a(FP_subtractor_13ccs_1_io_in_a),
    .io_in_b(FP_subtractor_13ccs_1_io_in_b),
    .io_out_s(FP_subtractor_13ccs_1_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_2 ( // @[FloatingPointDesigns.scala 2098:54]
    .clock(FP_subtractor_13ccs_2_clock),
    .reset(FP_subtractor_13ccs_2_reset),
    .io_in_a(FP_subtractor_13ccs_2_io_in_a),
    .io_in_b(FP_subtractor_13ccs_2_io_in_b),
    .io_out_s(FP_subtractor_13ccs_2_io_out_s)
  );
  assign io_out_s = {stage3_regs_r_1_1_8[31],FP_multiplier_10ccs_6_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2154:58]
  assign FP_multiplier_10ccs_clock = clock;
  assign FP_multiplier_10ccs_reset = reset;
  assign FP_multiplier_10ccs_io_in_a = {1'h0,result[30:0]}; // @[FloatingPointDesigns.scala 2034:48]
  assign FP_multiplier_10ccs_io_in_b = {1'h0,result[30:0]}; // @[FloatingPointDesigns.scala 2035:48]
  assign FP_multiplier_10ccs_1_clock = clock;
  assign FP_multiplier_10ccs_1_reset = reset;
  assign FP_multiplier_10ccs_1_io_in_a = FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2047:34]
  assign FP_multiplier_10ccs_1_io_in_b = {1'h0,stage1_regs_0_1_8[30:0]}; // @[FloatingPointDesigns.scala 2048:46]
  assign FP_multiplier_10ccs_2_clock = clock;
  assign FP_multiplier_10ccs_2_reset = reset;
  assign FP_multiplier_10ccs_2_io_in_a = {1'h0,stage3_regs_0_0_11[30:0]}; // @[FloatingPointDesigns.scala 2065:46]
  assign FP_multiplier_10ccs_2_io_in_b = FP_subtractor_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2066:34]
  assign FP_subtractor_13ccs_clock = clock;
  assign FP_subtractor_13ccs_reset = reset;
  assign FP_subtractor_13ccs_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1983:26 1984:16]
  assign FP_subtractor_13ccs_io_in_b = FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2057:31]
  assign multiplier4_clock = clock;
  assign multiplier4_reset = reset;
  assign multiplier4_io_in_a = {1'h0,FP_multiplier_10ccs_2_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2087:37]
  assign multiplier4_io_in_b = {1'h0,FP_multiplier_10ccs_2_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2088:37]
  assign FP_multiplier_10ccs_3_clock = clock;
  assign FP_multiplier_10ccs_3_reset = reset;
  assign FP_multiplier_10ccs_3_io_in_a = {1'h0,multiplier4_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2123:50]
  assign FP_multiplier_10ccs_3_io_in_b = {1'h0,transition_regs_8[30:0]}; // @[FloatingPointDesigns.scala 2124:50]
  assign FP_multiplier_10ccs_4_clock = clock;
  assign FP_multiplier_10ccs_4_reset = reset;
  assign FP_multiplier_10ccs_4_io_in_a = {1'h0,stage2_regs_r_0_0_11[30:0]}; // @[FloatingPointDesigns.scala 2145:48]
  assign FP_multiplier_10ccs_4_io_in_b = FP_subtractor_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2146:36]
  assign FP_multiplier_10ccs_5_clock = clock;
  assign FP_multiplier_10ccs_5_reset = reset;
  assign FP_multiplier_10ccs_5_io_in_a = {1'h0,FP_multiplier_10ccs_4_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2132:50]
  assign FP_multiplier_10ccs_5_io_in_b = {1'h0,stage3_regs_r_0_1_8[30:0]}; // @[FloatingPointDesigns.scala 2133:50]
  assign FP_multiplier_10ccs_6_clock = clock;
  assign FP_multiplier_10ccs_6_reset = reset;
  assign FP_multiplier_10ccs_6_io_in_a = {1'h0,stage2_regs_r_1_0_11[30:0]}; // @[FloatingPointDesigns.scala 2145:48]
  assign FP_multiplier_10ccs_6_io_in_b = FP_subtractor_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2146:36]
  assign FP_subtractor_13ccs_1_clock = clock;
  assign FP_subtractor_13ccs_1_reset = reset;
  assign FP_subtractor_13ccs_1_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 1985:19 1986:9]
  assign FP_subtractor_13ccs_1_io_in_b = FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2137:33]
  assign FP_subtractor_13ccs_2_clock = clock;
  assign FP_subtractor_13ccs_2_reset = reset;
  assign FP_subtractor_13ccs_2_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 1985:19 1986:9]
  assign FP_subtractor_13ccs_2_io_in_b = FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2137:33]
  always @(posedge clock) begin
    if (reset) begin // @[FloatingPointDesigns.scala 1999:22]
      x_n_0 <= 32'h0; // @[FloatingPointDesigns.scala 1999:22]
    end else begin
      x_n_0 <= result;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1999:22]
      x_n_1 <= 32'h0; // @[FloatingPointDesigns.scala 1999:22]
    end else begin
      x_n_1 <= stage1_regs_0_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1999:22]
      x_n_2 <= 32'h0; // @[FloatingPointDesigns.scala 1999:22]
    end else begin
      x_n_2 <= stage2_regs_0_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2000:22]
      a_2_0 <= 32'h0; // @[FloatingPointDesigns.scala 2000:22]
    end else begin
      a_2_0 <= _a_2_0_T_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2000:22]
      a_2_1 <= 32'h0; // @[FloatingPointDesigns.scala 2000:22]
    end else begin
      a_2_1 <= stage1_regs_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2000:22]
      a_2_2 <= 32'h0; // @[FloatingPointDesigns.scala 2000:22]
    end else begin
      a_2_2 <= stage2_regs_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2000:22]
      a_2_3 <= 32'h0; // @[FloatingPointDesigns.scala 2000:22]
    end else begin
      a_2_3 <= stage3_regs_0_1_11;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_0_0 <= x_n_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_0_1 <= stage1_regs_0_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_0_2 <= stage1_regs_0_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_0_3 <= stage1_regs_0_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_0_4 <= stage1_regs_0_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_0_5 <= stage1_regs_0_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_0_6 <= stage1_regs_0_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_0_7 <= stage1_regs_0_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_0_8 <= stage1_regs_0_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_1_0 <= a_2_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_1_1 <= stage1_regs_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_1_2 <= stage1_regs_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_1_3 <= stage1_regs_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_1_4 <= stage1_regs_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_1_5 <= stage1_regs_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_1_6 <= stage1_regs_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_1_7 <= stage1_regs_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:30]
      stage1_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2001:30]
    end else begin
      stage1_regs_0_1_8 <= stage1_regs_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_0_0 <= x_n_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_0_1 <= stage2_regs_0_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_0_2 <= stage2_regs_0_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_0_3 <= stage2_regs_0_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_0_4 <= stage2_regs_0_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_0_5 <= stage2_regs_0_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_0_6 <= stage2_regs_0_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_0_7 <= stage2_regs_0_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_0_8 <= stage2_regs_0_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_1_0 <= a_2_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_1_1 <= stage2_regs_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_1_2 <= stage2_regs_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_1_3 <= stage2_regs_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_1_4 <= stage2_regs_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_1_5 <= stage2_regs_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_1_6 <= stage2_regs_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_1_7 <= stage2_regs_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:30]
      stage2_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2002:30]
    end else begin
      stage2_regs_0_1_8 <= stage2_regs_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_0_0 <= x_n_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_0_1 <= stage3_regs_0_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_0_2 <= stage3_regs_0_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_0_3 <= stage3_regs_0_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_0_4 <= stage3_regs_0_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_0_5 <= stage3_regs_0_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_0_6 <= stage3_regs_0_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_0_7 <= stage3_regs_0_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_0_8 <= stage3_regs_0_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_0_9 <= stage3_regs_0_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_0_10 <= stage3_regs_0_0_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_0_11 <= stage3_regs_0_0_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_1_0 <= a_2_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_1_1 <= stage3_regs_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_1_2 <= stage3_regs_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_1_3 <= stage3_regs_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_1_4 <= stage3_regs_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_1_5 <= stage3_regs_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_1_6 <= stage3_regs_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_1_7 <= stage3_regs_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_1_8 <= stage3_regs_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_1_9 <= stage3_regs_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_1_10 <= stage3_regs_0_1_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage3_regs_0_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage3_regs_0_1_11 <= stage3_regs_0_1_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage4_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage4_regs_0_1_0 <= a_2_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage4_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage4_regs_0_1_1 <= stage4_regs_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage4_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage4_regs_0_1_2 <= stage4_regs_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage4_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage4_regs_0_1_3 <= stage4_regs_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage4_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage4_regs_0_1_4 <= stage4_regs_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage4_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage4_regs_0_1_5 <= stage4_regs_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage4_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage4_regs_0_1_6 <= stage4_regs_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage4_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage4_regs_0_1_7 <= stage4_regs_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage4_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage4_regs_0_1_8 <= stage4_regs_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2075:31]
      a_2_isr_to_r <= 32'h0; // @[FloatingPointDesigns.scala 2075:31]
    end else begin
      a_2_isr_to_r <= _a_2_isr_to_r_T_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2076:34]
      transition_regs_0 <= 32'h0; // @[FloatingPointDesigns.scala 2076:34]
    end else begin
      transition_regs_0 <= a_2_isr_to_r;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2076:34]
      transition_regs_1 <= 32'h0; // @[FloatingPointDesigns.scala 2076:34]
    end else begin
      transition_regs_1 <= transition_regs_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2076:34]
      transition_regs_2 <= 32'h0; // @[FloatingPointDesigns.scala 2076:34]
    end else begin
      transition_regs_2 <= transition_regs_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2076:34]
      transition_regs_3 <= 32'h0; // @[FloatingPointDesigns.scala 2076:34]
    end else begin
      transition_regs_3 <= transition_regs_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2076:34]
      transition_regs_4 <= 32'h0; // @[FloatingPointDesigns.scala 2076:34]
    end else begin
      transition_regs_4 <= transition_regs_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2076:34]
      transition_regs_5 <= 32'h0; // @[FloatingPointDesigns.scala 2076:34]
    end else begin
      transition_regs_5 <= transition_regs_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2076:34]
      transition_regs_6 <= 32'h0; // @[FloatingPointDesigns.scala 2076:34]
    end else begin
      transition_regs_6 <= transition_regs_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2076:34]
      transition_regs_7 <= 32'h0; // @[FloatingPointDesigns.scala 2076:34]
    end else begin
      transition_regs_7 <= transition_regs_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2076:34]
      transition_regs_8 <= 32'h0; // @[FloatingPointDesigns.scala 2076:34]
    end else begin
      transition_regs_8 <= transition_regs_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2092:24]
      x_n_r_0 <= 32'h0; // @[FloatingPointDesigns.scala 2092:24]
    end else begin
      x_n_r_0 <= _GEN_133;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2092:24]
      x_n_r_1 <= 32'h0; // @[FloatingPointDesigns.scala 2092:24]
    end else begin
      x_n_r_1 <= stage1_regs_r_0_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2092:24]
      x_n_r_3 <= 32'h0; // @[FloatingPointDesigns.scala 2092:24]
    end else begin
      x_n_r_3 <= _GEN_189;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2092:24]
      x_n_r_4 <= 32'h0; // @[FloatingPointDesigns.scala 2092:24]
    end else begin
      x_n_r_4 <= stage1_regs_r_1_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2093:24]
      a_2_r_0 <= 32'h0; // @[FloatingPointDesigns.scala 2093:24]
    end else begin
      a_2_r_0 <= transition_regs_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2093:24]
      a_2_r_1 <= 32'h0; // @[FloatingPointDesigns.scala 2093:24]
    end else begin
      a_2_r_1 <= stage1_regs_r_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2093:24]
      a_2_r_2 <= 32'h0; // @[FloatingPointDesigns.scala 2093:24]
    end else begin
      a_2_r_2 <= stage2_regs_r_0_1_11;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2093:24]
      a_2_r_3 <= 32'h0; // @[FloatingPointDesigns.scala 2093:24]
    end else begin
      a_2_r_3 <= stage3_regs_r_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2093:24]
      a_2_r_4 <= 32'h0; // @[FloatingPointDesigns.scala 2093:24]
    end else begin
      a_2_r_4 <= stage1_regs_r_1_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2093:24]
      a_2_r_5 <= 32'h0; // @[FloatingPointDesigns.scala 2093:24]
    end else begin
      a_2_r_5 <= stage2_regs_r_1_1_11;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_0_0 <= x_n_r_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_0_1 <= stage1_regs_r_0_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_0_2 <= stage1_regs_r_0_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_0_3 <= stage1_regs_r_0_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_0_4 <= stage1_regs_r_0_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_0_5 <= stage1_regs_r_0_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_0_6 <= stage1_regs_r_0_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_0_7 <= stage1_regs_r_0_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_0_8 <= stage1_regs_r_0_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_1_0 <= a_2_r_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_1_1 <= stage1_regs_r_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_1_2 <= stage1_regs_r_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_1_3 <= stage1_regs_r_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_1_4 <= stage1_regs_r_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_1_5 <= stage1_regs_r_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_1_6 <= stage1_regs_r_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_1_7 <= stage1_regs_r_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_0_1_8 <= stage1_regs_r_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_0_0 <= x_n_r_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_0_1 <= stage1_regs_r_1_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_0_2 <= stage1_regs_r_1_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_0_3 <= stage1_regs_r_1_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_0_4 <= stage1_regs_r_1_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_0_5 <= stage1_regs_r_1_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_0_6 <= stage1_regs_r_1_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_0_7 <= stage1_regs_r_1_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_0_8 <= stage1_regs_r_1_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_1_0 <= a_2_r_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_1_1 <= stage1_regs_r_1_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_1_2 <= stage1_regs_r_1_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_1_3 <= stage1_regs_r_1_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_1_4 <= stage1_regs_r_1_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_1_5 <= stage1_regs_r_1_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_1_6 <= stage1_regs_r_1_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_1_7 <= stage1_regs_r_1_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:32]
      stage1_regs_r_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2094:32]
    end else begin
      stage1_regs_r_1_1_8 <= stage1_regs_r_1_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_0_0 <= x_n_r_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_0_1 <= stage2_regs_r_0_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_0_2 <= stage2_regs_r_0_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_0_3 <= stage2_regs_r_0_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_0_4 <= stage2_regs_r_0_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_0_5 <= stage2_regs_r_0_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_0_6 <= stage2_regs_r_0_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_0_7 <= stage2_regs_r_0_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_0_8 <= stage2_regs_r_0_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_0_9 <= stage2_regs_r_0_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_0_10 <= stage2_regs_r_0_0_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_0_11 <= stage2_regs_r_0_0_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_1_0 <= a_2_r_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_1_1 <= stage2_regs_r_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_1_2 <= stage2_regs_r_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_1_3 <= stage2_regs_r_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_1_4 <= stage2_regs_r_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_1_5 <= stage2_regs_r_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_1_6 <= stage2_regs_r_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_1_7 <= stage2_regs_r_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_1_8 <= stage2_regs_r_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_1_9 <= stage2_regs_r_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_1_10 <= stage2_regs_r_0_1_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_0_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_0_1_11 <= stage2_regs_r_0_1_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_0_0 <= x_n_r_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_0_1 <= stage2_regs_r_1_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_0_2 <= stage2_regs_r_1_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_0_3 <= stage2_regs_r_1_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_0_4 <= stage2_regs_r_1_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_0_5 <= stage2_regs_r_1_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_0_6 <= stage2_regs_r_1_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_0_7 <= stage2_regs_r_1_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_0_8 <= stage2_regs_r_1_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_0_9 <= stage2_regs_r_1_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_0_10 <= stage2_regs_r_1_0_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_0_11 <= stage2_regs_r_1_0_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_1_0 <= a_2_r_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_1_1 <= stage2_regs_r_1_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_1_2 <= stage2_regs_r_1_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_1_3 <= stage2_regs_r_1_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_1_4 <= stage2_regs_r_1_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_1_5 <= stage2_regs_r_1_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_1_6 <= stage2_regs_r_1_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_1_7 <= stage2_regs_r_1_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_1_8 <= stage2_regs_r_1_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_1_9 <= stage2_regs_r_1_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_1_10 <= stage2_regs_r_1_1_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:32]
      stage2_regs_r_1_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2095:32]
    end else begin
      stage2_regs_r_1_1_11 <= stage2_regs_r_1_1_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_0_1_0 <= a_2_r_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_0_1_1 <= stage3_regs_r_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_0_1_2 <= stage3_regs_r_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_0_1_3 <= stage3_regs_r_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_0_1_4 <= stage3_regs_r_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_0_1_5 <= stage3_regs_r_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_0_1_6 <= stage3_regs_r_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_0_1_7 <= stage3_regs_r_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_0_1_8 <= stage3_regs_r_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_1_1_0 <= a_2_r_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_1_1_1 <= stage3_regs_r_1_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_1_1_2 <= stage3_regs_r_1_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_1_1_3 <= stage3_regs_r_1_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_1_1_4 <= stage3_regs_r_1_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_1_1_5 <= stage3_regs_r_1_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_1_1_6 <= stage3_regs_r_1_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_1_1_7 <= stage3_regs_r_1_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage3_regs_r_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage3_regs_r_1_1_8 <= stage3_regs_r_1_1_7;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  x_n_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  x_n_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  x_n_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  a_2_0 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  a_2_1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  a_2_2 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  a_2_3 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  stage1_regs_0_0_0 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  stage1_regs_0_0_1 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  stage1_regs_0_0_2 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  stage1_regs_0_0_3 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  stage1_regs_0_0_4 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  stage1_regs_0_0_5 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  stage1_regs_0_0_6 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  stage1_regs_0_0_7 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  stage1_regs_0_0_8 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  stage1_regs_0_1_0 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  stage1_regs_0_1_1 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  stage1_regs_0_1_2 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  stage1_regs_0_1_3 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  stage1_regs_0_1_4 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  stage1_regs_0_1_5 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  stage1_regs_0_1_6 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  stage1_regs_0_1_7 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  stage1_regs_0_1_8 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  stage2_regs_0_0_0 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  stage2_regs_0_0_1 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  stage2_regs_0_0_2 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  stage2_regs_0_0_3 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  stage2_regs_0_0_4 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  stage2_regs_0_0_5 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  stage2_regs_0_0_6 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  stage2_regs_0_0_7 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  stage2_regs_0_0_8 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  stage2_regs_0_1_0 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  stage2_regs_0_1_1 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  stage2_regs_0_1_2 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  stage2_regs_0_1_3 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  stage2_regs_0_1_4 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  stage2_regs_0_1_5 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  stage2_regs_0_1_6 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  stage2_regs_0_1_7 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  stage2_regs_0_1_8 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  stage3_regs_0_0_0 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  stage3_regs_0_0_1 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  stage3_regs_0_0_2 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  stage3_regs_0_0_3 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  stage3_regs_0_0_4 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  stage3_regs_0_0_5 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  stage3_regs_0_0_6 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  stage3_regs_0_0_7 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  stage3_regs_0_0_8 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  stage3_regs_0_0_9 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  stage3_regs_0_0_10 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  stage3_regs_0_0_11 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  stage3_regs_0_1_0 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  stage3_regs_0_1_1 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  stage3_regs_0_1_2 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  stage3_regs_0_1_3 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  stage3_regs_0_1_4 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  stage3_regs_0_1_5 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  stage3_regs_0_1_6 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  stage3_regs_0_1_7 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  stage3_regs_0_1_8 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  stage3_regs_0_1_9 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  stage3_regs_0_1_10 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  stage3_regs_0_1_11 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  stage4_regs_0_1_0 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  stage4_regs_0_1_1 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  stage4_regs_0_1_2 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  stage4_regs_0_1_3 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  stage4_regs_0_1_4 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  stage4_regs_0_1_5 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  stage4_regs_0_1_6 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  stage4_regs_0_1_7 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  stage4_regs_0_1_8 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  a_2_isr_to_r = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  transition_regs_0 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  transition_regs_1 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  transition_regs_2 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  transition_regs_3 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  transition_regs_4 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  transition_regs_5 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  transition_regs_6 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  transition_regs_7 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  transition_regs_8 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  x_n_r_0 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  x_n_r_1 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  x_n_r_3 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  x_n_r_4 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  a_2_r_0 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  a_2_r_1 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  a_2_r_2 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  a_2_r_3 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  a_2_r_4 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  a_2_r_5 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  stage1_regs_r_0_0_0 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  stage1_regs_r_0_0_1 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  stage1_regs_r_0_0_2 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  stage1_regs_r_0_0_3 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  stage1_regs_r_0_0_4 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  stage1_regs_r_0_0_5 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  stage1_regs_r_0_0_6 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  stage1_regs_r_0_0_7 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  stage1_regs_r_0_0_8 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  stage1_regs_r_0_1_0 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  stage1_regs_r_0_1_1 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  stage1_regs_r_0_1_2 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  stage1_regs_r_0_1_3 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  stage1_regs_r_0_1_4 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  stage1_regs_r_0_1_5 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  stage1_regs_r_0_1_6 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  stage1_regs_r_0_1_7 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  stage1_regs_r_0_1_8 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  stage1_regs_r_1_0_0 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  stage1_regs_r_1_0_1 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  stage1_regs_r_1_0_2 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  stage1_regs_r_1_0_3 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  stage1_regs_r_1_0_4 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  stage1_regs_r_1_0_5 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  stage1_regs_r_1_0_6 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  stage1_regs_r_1_0_7 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  stage1_regs_r_1_0_8 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  stage1_regs_r_1_1_0 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  stage1_regs_r_1_1_1 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  stage1_regs_r_1_1_2 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  stage1_regs_r_1_1_3 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  stage1_regs_r_1_1_4 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  stage1_regs_r_1_1_5 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  stage1_regs_r_1_1_6 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  stage1_regs_r_1_1_7 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  stage1_regs_r_1_1_8 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  stage2_regs_r_0_0_0 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  stage2_regs_r_0_0_1 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  stage2_regs_r_0_0_2 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  stage2_regs_r_0_0_3 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  stage2_regs_r_0_0_4 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  stage2_regs_r_0_0_5 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  stage2_regs_r_0_0_6 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  stage2_regs_r_0_0_7 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  stage2_regs_r_0_0_8 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  stage2_regs_r_0_0_9 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  stage2_regs_r_0_0_10 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  stage2_regs_r_0_0_11 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  stage2_regs_r_0_1_0 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  stage2_regs_r_0_1_1 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  stage2_regs_r_0_1_2 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  stage2_regs_r_0_1_3 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  stage2_regs_r_0_1_4 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  stage2_regs_r_0_1_5 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  stage2_regs_r_0_1_6 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  stage2_regs_r_0_1_7 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  stage2_regs_r_0_1_8 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  stage2_regs_r_0_1_9 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  stage2_regs_r_0_1_10 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  stage2_regs_r_0_1_11 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  stage2_regs_r_1_0_0 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  stage2_regs_r_1_0_1 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  stage2_regs_r_1_0_2 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  stage2_regs_r_1_0_3 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  stage2_regs_r_1_0_4 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  stage2_regs_r_1_0_5 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  stage2_regs_r_1_0_6 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  stage2_regs_r_1_0_7 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  stage2_regs_r_1_0_8 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  stage2_regs_r_1_0_9 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  stage2_regs_r_1_0_10 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  stage2_regs_r_1_0_11 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  stage2_regs_r_1_1_0 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  stage2_regs_r_1_1_1 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  stage2_regs_r_1_1_2 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  stage2_regs_r_1_1_3 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  stage2_regs_r_1_1_4 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  stage2_regs_r_1_1_5 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  stage2_regs_r_1_1_6 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  stage2_regs_r_1_1_7 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  stage2_regs_r_1_1_8 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  stage2_regs_r_1_1_9 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  stage2_regs_r_1_1_10 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  stage2_regs_r_1_1_11 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  stage3_regs_r_0_1_0 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  stage3_regs_r_0_1_1 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  stage3_regs_r_0_1_2 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  stage3_regs_r_0_1_3 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  stage3_regs_r_0_1_4 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  stage3_regs_r_0_1_5 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  stage3_regs_r_0_1_6 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  stage3_regs_r_0_1_7 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  stage3_regs_r_0_1_8 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  stage3_regs_r_1_1_0 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  stage3_regs_r_1_1_1 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  stage3_regs_r_1_1_2 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  stage3_regs_r_1_1_3 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  stage3_regs_r_1_1_4 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  stage3_regs_r_1_1_5 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  stage3_regs_r_1_1_6 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  stage3_regs_r_1_1_7 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  stage3_regs_r_1_1_8 = _RAND_197[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module hqr7(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  output [31:0] io_out_s
);
  wire  FP_multiplier_10ccs_clock; // @[FloatingPointDesigns.scala 2531:28]
  wire  FP_multiplier_10ccs_reset; // @[FloatingPointDesigns.scala 2531:28]
  wire [31:0] FP_multiplier_10ccs_io_in_a; // @[FloatingPointDesigns.scala 2531:28]
  wire [31:0] FP_multiplier_10ccs_io_in_b; // @[FloatingPointDesigns.scala 2531:28]
  wire [31:0] FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2531:28]
  wire  FP_reciprocal_newfpu_clock; // @[FloatingPointDesigns.scala 2532:28]
  wire  FP_reciprocal_newfpu_reset; // @[FloatingPointDesigns.scala 2532:28]
  wire [31:0] FP_reciprocal_newfpu_io_in_a; // @[FloatingPointDesigns.scala 2532:28]
  wire [31:0] FP_reciprocal_newfpu_io_out_s; // @[FloatingPointDesigns.scala 2532:28]
  FP_multiplier_10ccs FP_multiplier_10ccs ( // @[FloatingPointDesigns.scala 2531:28]
    .clock(FP_multiplier_10ccs_clock),
    .reset(FP_multiplier_10ccs_reset),
    .io_in_a(FP_multiplier_10ccs_io_in_a),
    .io_in_b(FP_multiplier_10ccs_io_in_b),
    .io_out_s(FP_multiplier_10ccs_io_out_s)
  );
  FP_reciprocal_newfpu FP_reciprocal_newfpu ( // @[FloatingPointDesigns.scala 2532:28]
    .clock(FP_reciprocal_newfpu_clock),
    .reset(FP_reciprocal_newfpu_reset),
    .io_in_a(FP_reciprocal_newfpu_io_in_a),
    .io_out_s(FP_reciprocal_newfpu_io_out_s)
  );
  assign io_out_s = FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2542:14]
  assign FP_multiplier_10ccs_clock = clock;
  assign FP_multiplier_10ccs_reset = reset;
  assign FP_multiplier_10ccs_io_in_a = 32'hc0000000; // @[FloatingPointDesigns.scala 2539:21]
  assign FP_multiplier_10ccs_io_in_b = FP_reciprocal_newfpu_io_out_s; // @[FloatingPointDesigns.scala 2540:21]
  assign FP_reciprocal_newfpu_clock = clock;
  assign FP_reciprocal_newfpu_reset = reset;
  assign FP_reciprocal_newfpu_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2537:21]
endmodule
module FPReg(
  input         clock,
  input         reset,
  input  [31:0] io_in,
  output [31:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_0; // @[FloatingPointDesigns.scala 2268:22]
  reg [31:0] reg_1; // @[FloatingPointDesigns.scala 2268:22]
  reg [31:0] reg_2; // @[FloatingPointDesigns.scala 2268:22]
  reg [31:0] reg_3; // @[FloatingPointDesigns.scala 2268:22]
  reg [31:0] reg_4; // @[FloatingPointDesigns.scala 2268:22]
  reg [31:0] reg_5; // @[FloatingPointDesigns.scala 2268:22]
  reg [31:0] reg_6; // @[FloatingPointDesigns.scala 2268:22]
  reg [31:0] reg_7; // @[FloatingPointDesigns.scala 2268:22]
  reg [31:0] reg_8; // @[FloatingPointDesigns.scala 2268:22]
  reg [31:0] reg_9; // @[FloatingPointDesigns.scala 2268:22]
  assign io_out = reg_9; // @[FloatingPointDesigns.scala 2274:12]
  always @(posedge clock) begin
    if (reset) begin // @[FloatingPointDesigns.scala 2268:22]
      reg_0 <= 32'h0; // @[FloatingPointDesigns.scala 2268:22]
    end else begin
      reg_0 <= io_in; // @[FloatingPointDesigns.scala 2270:14]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2268:22]
      reg_1 <= 32'h0; // @[FloatingPointDesigns.scala 2268:22]
    end else begin
      reg_1 <= reg_0; // @[FloatingPointDesigns.scala 2272:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2268:22]
      reg_2 <= 32'h0; // @[FloatingPointDesigns.scala 2268:22]
    end else begin
      reg_2 <= reg_1; // @[FloatingPointDesigns.scala 2272:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2268:22]
      reg_3 <= 32'h0; // @[FloatingPointDesigns.scala 2268:22]
    end else begin
      reg_3 <= reg_2; // @[FloatingPointDesigns.scala 2272:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2268:22]
      reg_4 <= 32'h0; // @[FloatingPointDesigns.scala 2268:22]
    end else begin
      reg_4 <= reg_3; // @[FloatingPointDesigns.scala 2272:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2268:22]
      reg_5 <= 32'h0; // @[FloatingPointDesigns.scala 2268:22]
    end else begin
      reg_5 <= reg_4; // @[FloatingPointDesigns.scala 2272:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2268:22]
      reg_6 <= 32'h0; // @[FloatingPointDesigns.scala 2268:22]
    end else begin
      reg_6 <= reg_5; // @[FloatingPointDesigns.scala 2272:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2268:22]
      reg_7 <= 32'h0; // @[FloatingPointDesigns.scala 2268:22]
    end else begin
      reg_7 <= reg_6; // @[FloatingPointDesigns.scala 2272:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2268:22]
      reg_8 <= 32'h0; // @[FloatingPointDesigns.scala 2268:22]
    end else begin
      reg_8 <= reg_7; // @[FloatingPointDesigns.scala 2272:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2268:22]
      reg_9 <= 32'h0; // @[FloatingPointDesigns.scala 2268:22]
    end else begin
      reg_9 <= reg_8; // @[FloatingPointDesigns.scala 2272:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_9 = _RAND_9[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module axpy_dp(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b_0,
  input  [31:0] io_in_b_1,
  input  [31:0] io_in_b_2,
  input  [31:0] io_in_b_3,
  input  [31:0] io_in_b_4,
  input  [31:0] io_in_b_5,
  input  [31:0] io_in_b_6,
  input  [31:0] io_in_b_7,
  input  [31:0] io_in_b_8,
  input  [31:0] io_in_b_9,
  input  [31:0] io_in_b_10,
  input  [31:0] io_in_b_11,
  input  [31:0] io_in_b_12,
  input  [31:0] io_in_b_13,
  input  [31:0] io_in_b_14,
  input  [31:0] io_in_b_15,
  input  [31:0] io_in_b_16,
  input  [31:0] io_in_b_17,
  input  [31:0] io_in_b_18,
  input  [31:0] io_in_b_19,
  input  [31:0] io_in_b_20,
  input  [31:0] io_in_b_21,
  input  [31:0] io_in_b_22,
  input  [31:0] io_in_b_23,
  input  [31:0] io_in_b_24,
  input  [31:0] io_in_b_25,
  input  [31:0] io_in_b_26,
  input  [31:0] io_in_b_27,
  input  [31:0] io_in_b_28,
  input  [31:0] io_in_b_29,
  input  [31:0] io_in_b_30,
  input  [31:0] io_in_b_31,
  input  [31:0] io_in_b_32,
  input  [31:0] io_in_b_33,
  input  [31:0] io_in_b_34,
  input  [31:0] io_in_b_35,
  input  [31:0] io_in_b_36,
  input  [31:0] io_in_b_37,
  input  [31:0] io_in_b_38,
  input  [31:0] io_in_b_39,
  input  [31:0] io_in_b_40,
  input  [31:0] io_in_b_41,
  input  [31:0] io_in_b_42,
  input  [31:0] io_in_b_43,
  input  [31:0] io_in_b_44,
  input  [31:0] io_in_b_45,
  input  [31:0] io_in_b_46,
  input  [31:0] io_in_b_47,
  input  [31:0] io_in_b_48,
  input  [31:0] io_in_b_49,
  input  [31:0] io_in_b_50,
  input  [31:0] io_in_b_51,
  input  [31:0] io_in_b_52,
  input  [31:0] io_in_b_53,
  input  [31:0] io_in_b_54,
  input  [31:0] io_in_b_55,
  input  [31:0] io_in_b_56,
  input  [31:0] io_in_b_57,
  input  [31:0] io_in_b_58,
  input  [31:0] io_in_b_59,
  input  [31:0] io_in_b_60,
  input  [31:0] io_in_b_61,
  input  [31:0] io_in_b_62,
  input  [31:0] io_in_b_63,
  input  [31:0] io_in_b_64,
  input  [31:0] io_in_b_65,
  input  [31:0] io_in_b_66,
  input  [31:0] io_in_b_67,
  input  [31:0] io_in_b_68,
  input  [31:0] io_in_b_69,
  input  [31:0] io_in_b_70,
  input  [31:0] io_in_b_71,
  input  [31:0] io_in_b_72,
  input  [31:0] io_in_b_73,
  input  [31:0] io_in_b_74,
  input  [31:0] io_in_b_75,
  input  [31:0] io_in_b_76,
  input  [31:0] io_in_b_77,
  input  [31:0] io_in_b_78,
  input  [31:0] io_in_b_79,
  input  [31:0] io_in_b_80,
  input  [31:0] io_in_b_81,
  input  [31:0] io_in_b_82,
  input  [31:0] io_in_b_83,
  input  [31:0] io_in_b_84,
  input  [31:0] io_in_b_85,
  input  [31:0] io_in_b_86,
  input  [31:0] io_in_b_87,
  input  [31:0] io_in_b_88,
  input  [31:0] io_in_b_89,
  input  [31:0] io_in_b_90,
  input  [31:0] io_in_b_91,
  input  [31:0] io_in_b_92,
  input  [31:0] io_in_b_93,
  input  [31:0] io_in_b_94,
  input  [31:0] io_in_b_95,
  input  [31:0] io_in_b_96,
  input  [31:0] io_in_b_97,
  input  [31:0] io_in_b_98,
  input  [31:0] io_in_b_99,
  input  [31:0] io_in_b_100,
  input  [31:0] io_in_b_101,
  input  [31:0] io_in_b_102,
  input  [31:0] io_in_b_103,
  input  [31:0] io_in_b_104,
  input  [31:0] io_in_b_105,
  input  [31:0] io_in_b_106,
  input  [31:0] io_in_b_107,
  input  [31:0] io_in_b_108,
  input  [31:0] io_in_b_109,
  input  [31:0] io_in_b_110,
  input  [31:0] io_in_b_111,
  input  [31:0] io_in_b_112,
  input  [31:0] io_in_b_113,
  input  [31:0] io_in_b_114,
  input  [31:0] io_in_b_115,
  input  [31:0] io_in_b_116,
  input  [31:0] io_in_b_117,
  input  [31:0] io_in_b_118,
  input  [31:0] io_in_b_119,
  input  [31:0] io_in_b_120,
  input  [31:0] io_in_b_121,
  input  [31:0] io_in_b_122,
  input  [31:0] io_in_b_123,
  input  [31:0] io_in_b_124,
  input  [31:0] io_in_b_125,
  input  [31:0] io_in_b_126,
  input  [31:0] io_in_b_127,
  input  [31:0] io_in_c_0,
  input  [31:0] io_in_c_1,
  input  [31:0] io_in_c_2,
  input  [31:0] io_in_c_3,
  input  [31:0] io_in_c_4,
  input  [31:0] io_in_c_5,
  input  [31:0] io_in_c_6,
  input  [31:0] io_in_c_7,
  input  [31:0] io_in_c_8,
  input  [31:0] io_in_c_9,
  input  [31:0] io_in_c_10,
  input  [31:0] io_in_c_11,
  input  [31:0] io_in_c_12,
  input  [31:0] io_in_c_13,
  input  [31:0] io_in_c_14,
  input  [31:0] io_in_c_15,
  input  [31:0] io_in_c_16,
  input  [31:0] io_in_c_17,
  input  [31:0] io_in_c_18,
  input  [31:0] io_in_c_19,
  input  [31:0] io_in_c_20,
  input  [31:0] io_in_c_21,
  input  [31:0] io_in_c_22,
  input  [31:0] io_in_c_23,
  input  [31:0] io_in_c_24,
  input  [31:0] io_in_c_25,
  input  [31:0] io_in_c_26,
  input  [31:0] io_in_c_27,
  input  [31:0] io_in_c_28,
  input  [31:0] io_in_c_29,
  input  [31:0] io_in_c_30,
  input  [31:0] io_in_c_31,
  input  [31:0] io_in_c_32,
  input  [31:0] io_in_c_33,
  input  [31:0] io_in_c_34,
  input  [31:0] io_in_c_35,
  input  [31:0] io_in_c_36,
  input  [31:0] io_in_c_37,
  input  [31:0] io_in_c_38,
  input  [31:0] io_in_c_39,
  input  [31:0] io_in_c_40,
  input  [31:0] io_in_c_41,
  input  [31:0] io_in_c_42,
  input  [31:0] io_in_c_43,
  input  [31:0] io_in_c_44,
  input  [31:0] io_in_c_45,
  input  [31:0] io_in_c_46,
  input  [31:0] io_in_c_47,
  input  [31:0] io_in_c_48,
  input  [31:0] io_in_c_49,
  input  [31:0] io_in_c_50,
  input  [31:0] io_in_c_51,
  input  [31:0] io_in_c_52,
  input  [31:0] io_in_c_53,
  input  [31:0] io_in_c_54,
  input  [31:0] io_in_c_55,
  input  [31:0] io_in_c_56,
  input  [31:0] io_in_c_57,
  input  [31:0] io_in_c_58,
  input  [31:0] io_in_c_59,
  input  [31:0] io_in_c_60,
  input  [31:0] io_in_c_61,
  input  [31:0] io_in_c_62,
  input  [31:0] io_in_c_63,
  input  [31:0] io_in_c_64,
  input  [31:0] io_in_c_65,
  input  [31:0] io_in_c_66,
  input  [31:0] io_in_c_67,
  input  [31:0] io_in_c_68,
  input  [31:0] io_in_c_69,
  input  [31:0] io_in_c_70,
  input  [31:0] io_in_c_71,
  input  [31:0] io_in_c_72,
  input  [31:0] io_in_c_73,
  input  [31:0] io_in_c_74,
  input  [31:0] io_in_c_75,
  input  [31:0] io_in_c_76,
  input  [31:0] io_in_c_77,
  input  [31:0] io_in_c_78,
  input  [31:0] io_in_c_79,
  input  [31:0] io_in_c_80,
  input  [31:0] io_in_c_81,
  input  [31:0] io_in_c_82,
  input  [31:0] io_in_c_83,
  input  [31:0] io_in_c_84,
  input  [31:0] io_in_c_85,
  input  [31:0] io_in_c_86,
  input  [31:0] io_in_c_87,
  input  [31:0] io_in_c_88,
  input  [31:0] io_in_c_89,
  input  [31:0] io_in_c_90,
  input  [31:0] io_in_c_91,
  input  [31:0] io_in_c_92,
  input  [31:0] io_in_c_93,
  input  [31:0] io_in_c_94,
  input  [31:0] io_in_c_95,
  input  [31:0] io_in_c_96,
  input  [31:0] io_in_c_97,
  input  [31:0] io_in_c_98,
  input  [31:0] io_in_c_99,
  input  [31:0] io_in_c_100,
  input  [31:0] io_in_c_101,
  input  [31:0] io_in_c_102,
  input  [31:0] io_in_c_103,
  input  [31:0] io_in_c_104,
  input  [31:0] io_in_c_105,
  input  [31:0] io_in_c_106,
  input  [31:0] io_in_c_107,
  input  [31:0] io_in_c_108,
  input  [31:0] io_in_c_109,
  input  [31:0] io_in_c_110,
  input  [31:0] io_in_c_111,
  input  [31:0] io_in_c_112,
  input  [31:0] io_in_c_113,
  input  [31:0] io_in_c_114,
  input  [31:0] io_in_c_115,
  input  [31:0] io_in_c_116,
  input  [31:0] io_in_c_117,
  input  [31:0] io_in_c_118,
  input  [31:0] io_in_c_119,
  input  [31:0] io_in_c_120,
  input  [31:0] io_in_c_121,
  input  [31:0] io_in_c_122,
  input  [31:0] io_in_c_123,
  input  [31:0] io_in_c_124,
  input  [31:0] io_in_c_125,
  input  [31:0] io_in_c_126,
  input  [31:0] io_in_c_127,
  output [31:0] io_out_s_0,
  output [31:0] io_out_s_1,
  output [31:0] io_out_s_2,
  output [31:0] io_out_s_3,
  output [31:0] io_out_s_4,
  output [31:0] io_out_s_5,
  output [31:0] io_out_s_6,
  output [31:0] io_out_s_7,
  output [31:0] io_out_s_8,
  output [31:0] io_out_s_9,
  output [31:0] io_out_s_10,
  output [31:0] io_out_s_11,
  output [31:0] io_out_s_12,
  output [31:0] io_out_s_13,
  output [31:0] io_out_s_14,
  output [31:0] io_out_s_15,
  output [31:0] io_out_s_16,
  output [31:0] io_out_s_17,
  output [31:0] io_out_s_18,
  output [31:0] io_out_s_19,
  output [31:0] io_out_s_20,
  output [31:0] io_out_s_21,
  output [31:0] io_out_s_22,
  output [31:0] io_out_s_23,
  output [31:0] io_out_s_24,
  output [31:0] io_out_s_25,
  output [31:0] io_out_s_26,
  output [31:0] io_out_s_27,
  output [31:0] io_out_s_28,
  output [31:0] io_out_s_29,
  output [31:0] io_out_s_30,
  output [31:0] io_out_s_31,
  output [31:0] io_out_s_32,
  output [31:0] io_out_s_33,
  output [31:0] io_out_s_34,
  output [31:0] io_out_s_35,
  output [31:0] io_out_s_36,
  output [31:0] io_out_s_37,
  output [31:0] io_out_s_38,
  output [31:0] io_out_s_39,
  output [31:0] io_out_s_40,
  output [31:0] io_out_s_41,
  output [31:0] io_out_s_42,
  output [31:0] io_out_s_43,
  output [31:0] io_out_s_44,
  output [31:0] io_out_s_45,
  output [31:0] io_out_s_46,
  output [31:0] io_out_s_47,
  output [31:0] io_out_s_48,
  output [31:0] io_out_s_49,
  output [31:0] io_out_s_50,
  output [31:0] io_out_s_51,
  output [31:0] io_out_s_52,
  output [31:0] io_out_s_53,
  output [31:0] io_out_s_54,
  output [31:0] io_out_s_55,
  output [31:0] io_out_s_56,
  output [31:0] io_out_s_57,
  output [31:0] io_out_s_58,
  output [31:0] io_out_s_59,
  output [31:0] io_out_s_60,
  output [31:0] io_out_s_61,
  output [31:0] io_out_s_62,
  output [31:0] io_out_s_63,
  output [31:0] io_out_s_64,
  output [31:0] io_out_s_65,
  output [31:0] io_out_s_66,
  output [31:0] io_out_s_67,
  output [31:0] io_out_s_68,
  output [31:0] io_out_s_69,
  output [31:0] io_out_s_70,
  output [31:0] io_out_s_71,
  output [31:0] io_out_s_72,
  output [31:0] io_out_s_73,
  output [31:0] io_out_s_74,
  output [31:0] io_out_s_75,
  output [31:0] io_out_s_76,
  output [31:0] io_out_s_77,
  output [31:0] io_out_s_78,
  output [31:0] io_out_s_79,
  output [31:0] io_out_s_80,
  output [31:0] io_out_s_81,
  output [31:0] io_out_s_82,
  output [31:0] io_out_s_83,
  output [31:0] io_out_s_84,
  output [31:0] io_out_s_85,
  output [31:0] io_out_s_86,
  output [31:0] io_out_s_87,
  output [31:0] io_out_s_88,
  output [31:0] io_out_s_89,
  output [31:0] io_out_s_90,
  output [31:0] io_out_s_91,
  output [31:0] io_out_s_92,
  output [31:0] io_out_s_93,
  output [31:0] io_out_s_94,
  output [31:0] io_out_s_95,
  output [31:0] io_out_s_96,
  output [31:0] io_out_s_97,
  output [31:0] io_out_s_98,
  output [31:0] io_out_s_99,
  output [31:0] io_out_s_100,
  output [31:0] io_out_s_101,
  output [31:0] io_out_s_102,
  output [31:0] io_out_s_103,
  output [31:0] io_out_s_104,
  output [31:0] io_out_s_105,
  output [31:0] io_out_s_106,
  output [31:0] io_out_s_107,
  output [31:0] io_out_s_108,
  output [31:0] io_out_s_109,
  output [31:0] io_out_s_110,
  output [31:0] io_out_s_111,
  output [31:0] io_out_s_112,
  output [31:0] io_out_s_113,
  output [31:0] io_out_s_114,
  output [31:0] io_out_s_115,
  output [31:0] io_out_s_116,
  output [31:0] io_out_s_117,
  output [31:0] io_out_s_118,
  output [31:0] io_out_s_119,
  output [31:0] io_out_s_120,
  output [31:0] io_out_s_121,
  output [31:0] io_out_s_122,
  output [31:0] io_out_s_123,
  output [31:0] io_out_s_124,
  output [31:0] io_out_s_125,
  output [31:0] io_out_s_126,
  output [31:0] io_out_s_127
);
  wire  FP_multiplier_10ccs_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_1_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_1_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_1_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_1_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_2_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_2_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_2_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_2_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_3_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_3_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_3_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_3_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_4_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_4_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_4_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_4_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_5_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_5_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_5_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_5_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_6_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_6_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_6_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_6_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_7_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_7_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_7_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_7_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_8_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_8_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_8_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_8_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_9_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_9_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_9_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_9_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_10_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_10_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_10_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_10_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_11_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_11_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_11_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_11_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_12_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_12_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_12_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_12_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_13_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_13_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_13_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_13_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_14_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_14_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_14_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_14_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_15_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_15_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_15_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_15_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_16_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_16_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_16_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_16_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_17_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_17_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_17_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_17_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_18_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_18_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_18_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_18_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_19_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_19_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_19_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_19_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_20_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_20_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_20_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_20_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_21_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_21_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_21_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_21_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_22_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_22_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_22_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_22_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_23_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_23_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_23_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_23_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_24_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_24_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_24_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_24_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_25_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_25_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_25_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_25_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_26_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_26_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_26_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_26_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_27_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_27_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_27_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_27_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_28_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_28_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_28_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_28_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_29_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_29_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_29_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_29_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_30_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_30_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_30_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_30_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_31_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_31_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_31_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_31_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_32_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_32_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_32_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_32_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_33_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_33_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_33_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_33_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_34_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_34_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_34_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_34_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_35_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_35_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_35_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_35_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_36_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_36_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_36_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_36_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_37_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_37_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_37_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_37_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_38_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_38_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_38_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_38_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_39_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_39_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_39_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_39_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_40_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_40_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_40_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_40_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_41_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_41_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_41_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_41_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_42_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_42_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_42_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_42_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_43_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_43_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_43_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_43_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_44_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_44_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_44_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_44_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_45_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_45_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_45_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_45_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_46_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_46_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_46_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_46_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_47_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_47_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_47_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_47_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_47_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_48_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_48_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_48_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_48_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_49_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_49_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_49_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_49_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_50_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_50_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_50_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_50_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_51_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_51_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_51_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_51_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_52_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_52_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_52_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_52_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_53_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_53_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_53_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_53_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_54_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_54_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_54_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_54_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_55_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_55_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_55_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_55_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_56_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_56_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_56_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_56_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_57_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_57_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_57_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_57_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_58_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_58_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_58_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_58_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_59_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_59_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_59_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_59_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_60_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_60_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_60_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_60_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_61_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_61_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_61_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_61_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_62_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_62_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_62_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_62_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_63_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_63_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_63_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_63_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_63_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_64_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_64_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_64_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_64_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_64_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_65_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_65_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_65_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_65_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_65_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_66_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_66_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_66_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_66_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_66_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_67_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_67_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_67_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_67_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_67_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_68_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_68_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_68_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_68_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_68_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_69_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_69_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_69_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_69_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_69_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_70_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_70_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_70_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_70_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_70_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_71_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_71_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_71_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_71_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_71_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_72_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_72_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_72_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_72_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_72_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_73_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_73_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_73_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_73_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_73_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_74_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_74_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_74_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_74_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_74_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_75_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_75_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_75_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_75_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_75_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_76_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_76_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_76_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_76_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_76_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_77_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_77_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_77_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_77_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_77_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_78_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_78_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_78_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_78_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_78_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_79_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_79_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_79_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_79_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_79_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_80_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_80_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_80_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_80_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_80_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_81_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_81_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_81_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_81_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_81_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_82_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_82_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_82_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_82_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_82_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_83_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_83_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_83_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_83_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_83_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_84_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_84_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_84_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_84_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_84_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_85_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_85_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_85_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_85_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_85_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_86_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_86_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_86_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_86_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_86_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_87_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_87_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_87_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_87_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_87_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_88_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_88_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_88_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_88_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_88_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_89_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_89_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_89_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_89_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_89_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_90_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_90_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_90_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_90_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_90_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_91_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_91_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_91_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_91_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_91_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_92_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_92_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_92_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_92_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_92_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_93_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_93_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_93_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_93_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_93_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_94_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_94_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_94_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_94_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_94_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_95_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_95_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_95_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_95_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_95_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_96_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_96_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_96_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_96_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_96_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_97_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_97_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_97_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_97_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_97_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_98_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_98_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_98_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_98_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_98_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_99_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_99_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_99_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_99_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_99_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_100_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_100_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_100_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_100_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_100_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_101_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_101_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_101_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_101_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_101_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_102_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_102_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_102_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_102_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_102_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_103_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_103_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_103_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_103_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_103_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_104_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_104_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_104_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_104_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_104_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_105_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_105_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_105_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_105_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_105_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_106_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_106_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_106_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_106_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_106_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_107_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_107_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_107_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_107_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_107_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_108_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_108_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_108_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_108_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_108_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_109_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_109_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_109_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_109_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_109_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_110_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_110_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_110_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_110_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_110_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_111_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_111_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_111_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_111_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_111_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_112_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_112_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_112_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_112_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_112_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_113_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_113_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_113_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_113_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_113_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_114_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_114_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_114_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_114_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_114_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_115_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_115_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_115_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_115_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_115_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_116_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_116_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_116_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_116_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_116_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_117_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_117_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_117_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_117_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_117_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_118_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_118_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_118_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_118_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_118_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_119_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_119_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_119_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_119_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_119_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_120_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_120_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_120_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_120_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_120_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_121_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_121_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_121_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_121_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_121_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_122_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_122_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_122_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_122_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_122_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_123_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_123_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_123_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_123_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_123_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_124_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_124_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_124_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_124_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_124_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_125_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_125_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_125_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_125_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_125_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_126_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_126_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_126_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_126_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_126_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_127_clock; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_multiplier_10ccs_127_reset; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_127_io_in_a; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_127_io_in_b; // @[FloatingPointDesigns.scala 2483:28]
  wire [31:0] FP_multiplier_10ccs_127_io_out_s; // @[FloatingPointDesigns.scala 2483:28]
  wire  FP_adder_13ccs_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_1_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_1_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_1_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_1_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_2_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_2_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_2_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_2_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_3_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_3_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_3_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_3_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_4_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_4_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_4_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_4_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_5_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_5_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_5_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_5_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_6_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_6_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_6_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_6_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_7_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_7_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_7_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_7_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_8_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_8_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_8_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_8_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_9_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_9_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_9_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_9_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_10_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_10_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_10_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_10_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_11_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_11_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_11_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_11_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_12_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_12_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_12_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_12_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_13_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_13_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_13_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_13_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_14_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_14_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_14_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_14_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_15_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_15_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_15_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_15_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_16_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_16_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_16_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_16_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_17_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_17_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_17_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_17_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_18_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_18_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_18_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_18_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_19_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_19_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_19_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_19_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_20_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_20_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_20_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_20_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_21_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_21_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_21_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_21_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_22_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_22_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_22_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_22_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_23_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_23_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_23_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_23_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_24_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_24_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_24_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_24_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_25_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_25_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_25_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_25_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_26_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_26_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_26_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_26_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_27_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_27_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_27_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_27_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_28_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_28_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_28_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_28_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_29_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_29_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_29_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_29_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_30_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_30_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_30_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_30_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_31_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_31_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_31_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_31_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_32_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_32_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_32_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_32_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_33_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_33_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_33_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_33_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_34_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_34_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_34_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_34_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_35_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_35_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_35_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_35_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_36_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_36_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_36_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_36_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_37_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_37_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_37_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_37_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_38_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_38_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_38_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_38_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_39_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_39_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_39_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_39_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_40_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_40_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_40_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_40_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_41_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_41_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_41_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_41_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_42_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_42_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_42_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_42_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_43_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_43_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_43_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_43_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_44_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_44_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_44_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_44_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_45_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_45_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_45_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_45_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_46_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_46_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_46_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_46_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_47_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_47_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_47_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_47_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_47_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_48_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_48_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_48_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_48_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_49_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_49_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_49_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_49_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_50_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_50_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_50_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_50_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_51_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_51_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_51_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_51_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_52_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_52_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_52_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_52_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_53_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_53_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_53_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_53_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_54_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_54_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_54_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_54_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_55_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_55_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_55_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_55_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_56_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_56_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_56_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_56_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_57_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_57_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_57_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_57_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_58_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_58_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_58_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_58_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_59_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_59_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_59_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_59_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_60_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_60_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_60_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_60_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_61_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_61_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_61_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_61_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_62_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_62_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_62_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_62_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_63_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_63_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_63_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_63_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_63_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_64_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_64_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_64_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_64_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_64_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_65_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_65_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_65_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_65_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_65_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_66_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_66_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_66_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_66_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_66_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_67_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_67_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_67_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_67_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_67_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_68_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_68_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_68_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_68_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_68_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_69_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_69_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_69_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_69_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_69_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_70_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_70_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_70_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_70_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_70_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_71_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_71_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_71_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_71_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_71_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_72_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_72_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_72_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_72_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_72_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_73_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_73_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_73_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_73_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_73_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_74_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_74_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_74_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_74_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_74_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_75_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_75_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_75_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_75_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_75_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_76_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_76_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_76_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_76_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_76_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_77_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_77_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_77_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_77_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_77_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_78_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_78_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_78_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_78_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_78_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_79_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_79_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_79_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_79_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_79_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_80_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_80_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_80_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_80_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_80_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_81_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_81_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_81_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_81_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_81_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_82_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_82_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_82_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_82_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_82_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_83_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_83_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_83_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_83_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_83_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_84_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_84_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_84_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_84_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_84_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_85_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_85_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_85_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_85_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_85_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_86_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_86_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_86_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_86_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_86_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_87_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_87_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_87_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_87_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_87_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_88_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_88_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_88_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_88_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_88_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_89_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_89_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_89_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_89_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_89_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_90_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_90_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_90_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_90_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_90_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_91_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_91_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_91_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_91_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_91_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_92_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_92_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_92_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_92_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_92_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_93_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_93_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_93_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_93_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_93_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_94_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_94_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_94_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_94_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_94_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_95_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_95_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_95_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_95_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_95_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_96_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_96_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_96_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_96_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_96_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_97_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_97_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_97_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_97_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_97_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_98_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_98_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_98_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_98_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_98_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_99_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_99_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_99_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_99_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_99_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_100_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_100_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_100_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_100_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_100_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_101_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_101_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_101_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_101_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_101_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_102_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_102_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_102_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_102_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_102_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_103_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_103_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_103_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_103_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_103_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_104_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_104_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_104_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_104_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_104_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_105_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_105_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_105_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_105_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_105_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_106_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_106_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_106_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_106_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_106_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_107_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_107_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_107_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_107_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_107_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_108_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_108_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_108_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_108_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_108_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_109_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_109_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_109_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_109_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_109_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_110_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_110_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_110_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_110_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_110_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_111_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_111_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_111_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_111_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_111_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_112_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_112_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_112_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_112_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_112_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_113_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_113_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_113_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_113_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_113_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_114_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_114_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_114_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_114_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_114_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_115_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_115_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_115_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_115_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_115_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_116_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_116_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_116_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_116_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_116_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_117_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_117_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_117_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_117_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_117_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_118_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_118_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_118_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_118_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_118_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_119_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_119_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_119_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_119_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_119_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_120_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_120_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_120_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_120_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_120_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_121_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_121_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_121_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_121_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_121_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_122_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_122_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_122_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_122_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_122_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_123_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_123_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_123_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_123_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_123_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_124_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_124_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_124_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_124_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_124_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_125_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_125_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_125_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_125_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_125_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_126_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_126_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_126_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_126_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_126_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_127_clock; // @[FloatingPointDesigns.scala 2488:25]
  wire  FP_adder_13ccs_127_reset; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_127_io_in_a; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_127_io_in_b; // @[FloatingPointDesigns.scala 2488:25]
  wire [31:0] FP_adder_13ccs_127_io_out_s; // @[FloatingPointDesigns.scala 2488:25]
  wire  FPReg_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_1_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_1_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_1_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_1_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_2_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_2_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_2_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_2_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_3_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_3_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_3_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_3_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_4_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_4_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_4_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_4_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_5_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_5_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_5_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_5_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_6_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_6_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_6_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_6_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_7_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_7_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_7_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_7_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_8_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_8_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_8_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_8_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_9_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_9_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_9_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_9_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_10_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_10_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_10_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_10_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_11_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_11_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_11_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_11_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_12_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_12_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_12_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_12_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_13_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_13_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_13_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_13_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_14_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_14_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_14_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_14_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_15_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_15_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_15_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_15_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_16_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_16_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_16_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_16_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_17_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_17_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_17_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_17_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_18_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_18_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_18_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_18_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_19_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_19_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_19_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_19_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_20_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_20_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_20_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_20_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_21_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_21_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_21_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_21_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_22_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_22_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_22_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_22_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_23_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_23_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_23_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_23_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_24_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_24_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_24_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_24_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_25_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_25_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_25_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_25_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_26_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_26_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_26_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_26_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_27_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_27_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_27_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_27_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_28_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_28_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_28_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_28_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_29_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_29_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_29_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_29_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_30_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_30_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_30_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_30_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_31_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_31_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_31_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_31_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_32_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_32_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_32_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_32_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_33_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_33_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_33_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_33_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_34_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_34_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_34_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_34_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_35_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_35_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_35_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_35_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_36_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_36_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_36_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_36_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_37_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_37_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_37_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_37_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_38_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_38_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_38_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_38_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_39_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_39_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_39_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_39_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_40_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_40_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_40_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_40_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_41_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_41_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_41_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_41_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_42_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_42_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_42_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_42_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_43_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_43_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_43_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_43_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_44_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_44_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_44_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_44_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_45_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_45_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_45_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_45_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_46_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_46_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_46_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_46_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_47_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_47_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_47_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_47_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_48_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_48_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_48_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_48_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_49_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_49_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_49_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_49_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_50_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_50_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_50_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_50_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_51_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_51_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_51_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_51_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_52_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_52_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_52_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_52_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_53_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_53_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_53_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_53_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_54_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_54_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_54_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_54_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_55_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_55_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_55_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_55_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_56_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_56_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_56_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_56_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_57_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_57_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_57_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_57_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_58_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_58_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_58_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_58_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_59_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_59_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_59_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_59_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_60_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_60_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_60_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_60_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_61_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_61_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_61_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_61_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_62_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_62_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_62_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_62_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_63_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_63_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_63_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_63_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_64_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_64_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_64_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_64_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_65_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_65_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_65_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_65_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_66_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_66_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_66_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_66_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_67_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_67_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_67_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_67_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_68_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_68_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_68_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_68_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_69_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_69_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_69_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_69_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_70_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_70_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_70_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_70_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_71_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_71_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_71_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_71_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_72_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_72_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_72_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_72_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_73_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_73_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_73_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_73_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_74_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_74_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_74_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_74_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_75_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_75_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_75_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_75_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_76_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_76_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_76_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_76_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_77_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_77_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_77_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_77_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_78_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_78_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_78_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_78_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_79_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_79_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_79_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_79_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_80_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_80_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_80_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_80_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_81_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_81_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_81_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_81_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_82_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_82_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_82_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_82_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_83_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_83_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_83_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_83_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_84_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_84_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_84_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_84_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_85_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_85_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_85_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_85_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_86_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_86_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_86_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_86_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_87_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_87_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_87_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_87_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_88_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_88_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_88_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_88_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_89_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_89_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_89_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_89_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_90_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_90_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_90_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_90_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_91_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_91_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_91_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_91_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_92_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_92_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_92_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_92_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_93_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_93_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_93_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_93_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_94_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_94_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_94_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_94_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_95_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_95_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_95_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_95_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_96_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_96_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_96_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_96_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_97_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_97_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_97_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_97_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_98_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_98_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_98_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_98_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_99_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_99_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_99_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_99_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_100_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_100_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_100_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_100_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_101_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_101_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_101_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_101_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_102_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_102_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_102_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_102_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_103_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_103_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_103_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_103_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_104_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_104_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_104_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_104_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_105_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_105_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_105_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_105_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_106_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_106_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_106_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_106_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_107_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_107_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_107_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_107_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_108_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_108_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_108_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_108_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_109_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_109_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_109_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_109_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_110_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_110_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_110_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_110_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_111_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_111_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_111_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_111_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_112_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_112_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_112_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_112_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_113_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_113_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_113_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_113_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_114_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_114_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_114_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_114_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_115_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_115_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_115_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_115_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_116_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_116_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_116_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_116_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_117_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_117_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_117_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_117_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_118_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_118_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_118_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_118_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_119_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_119_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_119_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_119_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_120_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_120_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_120_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_120_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_121_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_121_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_121_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_121_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_122_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_122_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_122_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_122_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_123_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_123_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_123_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_123_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_124_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_124_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_124_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_124_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_125_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_125_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_125_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_125_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_126_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_126_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_126_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_126_io_out; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_127_clock; // @[FloatingPointDesigns.scala 2492:48]
  wire  FPReg_127_reset; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_127_io_in; // @[FloatingPointDesigns.scala 2492:48]
  wire [31:0] FPReg_127_io_out; // @[FloatingPointDesigns.scala 2492:48]
  FP_multiplier_10ccs FP_multiplier_10ccs ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_clock),
    .reset(FP_multiplier_10ccs_reset),
    .io_in_a(FP_multiplier_10ccs_io_in_a),
    .io_in_b(FP_multiplier_10ccs_io_in_b),
    .io_out_s(FP_multiplier_10ccs_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_1 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_1_clock),
    .reset(FP_multiplier_10ccs_1_reset),
    .io_in_a(FP_multiplier_10ccs_1_io_in_a),
    .io_in_b(FP_multiplier_10ccs_1_io_in_b),
    .io_out_s(FP_multiplier_10ccs_1_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_2 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_2_clock),
    .reset(FP_multiplier_10ccs_2_reset),
    .io_in_a(FP_multiplier_10ccs_2_io_in_a),
    .io_in_b(FP_multiplier_10ccs_2_io_in_b),
    .io_out_s(FP_multiplier_10ccs_2_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_3 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_3_clock),
    .reset(FP_multiplier_10ccs_3_reset),
    .io_in_a(FP_multiplier_10ccs_3_io_in_a),
    .io_in_b(FP_multiplier_10ccs_3_io_in_b),
    .io_out_s(FP_multiplier_10ccs_3_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_4 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_4_clock),
    .reset(FP_multiplier_10ccs_4_reset),
    .io_in_a(FP_multiplier_10ccs_4_io_in_a),
    .io_in_b(FP_multiplier_10ccs_4_io_in_b),
    .io_out_s(FP_multiplier_10ccs_4_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_5 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_5_clock),
    .reset(FP_multiplier_10ccs_5_reset),
    .io_in_a(FP_multiplier_10ccs_5_io_in_a),
    .io_in_b(FP_multiplier_10ccs_5_io_in_b),
    .io_out_s(FP_multiplier_10ccs_5_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_6 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_6_clock),
    .reset(FP_multiplier_10ccs_6_reset),
    .io_in_a(FP_multiplier_10ccs_6_io_in_a),
    .io_in_b(FP_multiplier_10ccs_6_io_in_b),
    .io_out_s(FP_multiplier_10ccs_6_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_7 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_7_clock),
    .reset(FP_multiplier_10ccs_7_reset),
    .io_in_a(FP_multiplier_10ccs_7_io_in_a),
    .io_in_b(FP_multiplier_10ccs_7_io_in_b),
    .io_out_s(FP_multiplier_10ccs_7_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_8 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_8_clock),
    .reset(FP_multiplier_10ccs_8_reset),
    .io_in_a(FP_multiplier_10ccs_8_io_in_a),
    .io_in_b(FP_multiplier_10ccs_8_io_in_b),
    .io_out_s(FP_multiplier_10ccs_8_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_9 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_9_clock),
    .reset(FP_multiplier_10ccs_9_reset),
    .io_in_a(FP_multiplier_10ccs_9_io_in_a),
    .io_in_b(FP_multiplier_10ccs_9_io_in_b),
    .io_out_s(FP_multiplier_10ccs_9_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_10 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_10_clock),
    .reset(FP_multiplier_10ccs_10_reset),
    .io_in_a(FP_multiplier_10ccs_10_io_in_a),
    .io_in_b(FP_multiplier_10ccs_10_io_in_b),
    .io_out_s(FP_multiplier_10ccs_10_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_11 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_11_clock),
    .reset(FP_multiplier_10ccs_11_reset),
    .io_in_a(FP_multiplier_10ccs_11_io_in_a),
    .io_in_b(FP_multiplier_10ccs_11_io_in_b),
    .io_out_s(FP_multiplier_10ccs_11_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_12 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_12_clock),
    .reset(FP_multiplier_10ccs_12_reset),
    .io_in_a(FP_multiplier_10ccs_12_io_in_a),
    .io_in_b(FP_multiplier_10ccs_12_io_in_b),
    .io_out_s(FP_multiplier_10ccs_12_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_13 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_13_clock),
    .reset(FP_multiplier_10ccs_13_reset),
    .io_in_a(FP_multiplier_10ccs_13_io_in_a),
    .io_in_b(FP_multiplier_10ccs_13_io_in_b),
    .io_out_s(FP_multiplier_10ccs_13_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_14 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_14_clock),
    .reset(FP_multiplier_10ccs_14_reset),
    .io_in_a(FP_multiplier_10ccs_14_io_in_a),
    .io_in_b(FP_multiplier_10ccs_14_io_in_b),
    .io_out_s(FP_multiplier_10ccs_14_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_15 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_15_clock),
    .reset(FP_multiplier_10ccs_15_reset),
    .io_in_a(FP_multiplier_10ccs_15_io_in_a),
    .io_in_b(FP_multiplier_10ccs_15_io_in_b),
    .io_out_s(FP_multiplier_10ccs_15_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_16 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_16_clock),
    .reset(FP_multiplier_10ccs_16_reset),
    .io_in_a(FP_multiplier_10ccs_16_io_in_a),
    .io_in_b(FP_multiplier_10ccs_16_io_in_b),
    .io_out_s(FP_multiplier_10ccs_16_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_17 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_17_clock),
    .reset(FP_multiplier_10ccs_17_reset),
    .io_in_a(FP_multiplier_10ccs_17_io_in_a),
    .io_in_b(FP_multiplier_10ccs_17_io_in_b),
    .io_out_s(FP_multiplier_10ccs_17_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_18 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_18_clock),
    .reset(FP_multiplier_10ccs_18_reset),
    .io_in_a(FP_multiplier_10ccs_18_io_in_a),
    .io_in_b(FP_multiplier_10ccs_18_io_in_b),
    .io_out_s(FP_multiplier_10ccs_18_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_19 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_19_clock),
    .reset(FP_multiplier_10ccs_19_reset),
    .io_in_a(FP_multiplier_10ccs_19_io_in_a),
    .io_in_b(FP_multiplier_10ccs_19_io_in_b),
    .io_out_s(FP_multiplier_10ccs_19_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_20 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_20_clock),
    .reset(FP_multiplier_10ccs_20_reset),
    .io_in_a(FP_multiplier_10ccs_20_io_in_a),
    .io_in_b(FP_multiplier_10ccs_20_io_in_b),
    .io_out_s(FP_multiplier_10ccs_20_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_21 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_21_clock),
    .reset(FP_multiplier_10ccs_21_reset),
    .io_in_a(FP_multiplier_10ccs_21_io_in_a),
    .io_in_b(FP_multiplier_10ccs_21_io_in_b),
    .io_out_s(FP_multiplier_10ccs_21_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_22 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_22_clock),
    .reset(FP_multiplier_10ccs_22_reset),
    .io_in_a(FP_multiplier_10ccs_22_io_in_a),
    .io_in_b(FP_multiplier_10ccs_22_io_in_b),
    .io_out_s(FP_multiplier_10ccs_22_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_23 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_23_clock),
    .reset(FP_multiplier_10ccs_23_reset),
    .io_in_a(FP_multiplier_10ccs_23_io_in_a),
    .io_in_b(FP_multiplier_10ccs_23_io_in_b),
    .io_out_s(FP_multiplier_10ccs_23_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_24 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_24_clock),
    .reset(FP_multiplier_10ccs_24_reset),
    .io_in_a(FP_multiplier_10ccs_24_io_in_a),
    .io_in_b(FP_multiplier_10ccs_24_io_in_b),
    .io_out_s(FP_multiplier_10ccs_24_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_25 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_25_clock),
    .reset(FP_multiplier_10ccs_25_reset),
    .io_in_a(FP_multiplier_10ccs_25_io_in_a),
    .io_in_b(FP_multiplier_10ccs_25_io_in_b),
    .io_out_s(FP_multiplier_10ccs_25_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_26 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_26_clock),
    .reset(FP_multiplier_10ccs_26_reset),
    .io_in_a(FP_multiplier_10ccs_26_io_in_a),
    .io_in_b(FP_multiplier_10ccs_26_io_in_b),
    .io_out_s(FP_multiplier_10ccs_26_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_27 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_27_clock),
    .reset(FP_multiplier_10ccs_27_reset),
    .io_in_a(FP_multiplier_10ccs_27_io_in_a),
    .io_in_b(FP_multiplier_10ccs_27_io_in_b),
    .io_out_s(FP_multiplier_10ccs_27_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_28 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_28_clock),
    .reset(FP_multiplier_10ccs_28_reset),
    .io_in_a(FP_multiplier_10ccs_28_io_in_a),
    .io_in_b(FP_multiplier_10ccs_28_io_in_b),
    .io_out_s(FP_multiplier_10ccs_28_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_29 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_29_clock),
    .reset(FP_multiplier_10ccs_29_reset),
    .io_in_a(FP_multiplier_10ccs_29_io_in_a),
    .io_in_b(FP_multiplier_10ccs_29_io_in_b),
    .io_out_s(FP_multiplier_10ccs_29_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_30 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_30_clock),
    .reset(FP_multiplier_10ccs_30_reset),
    .io_in_a(FP_multiplier_10ccs_30_io_in_a),
    .io_in_b(FP_multiplier_10ccs_30_io_in_b),
    .io_out_s(FP_multiplier_10ccs_30_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_31 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_31_clock),
    .reset(FP_multiplier_10ccs_31_reset),
    .io_in_a(FP_multiplier_10ccs_31_io_in_a),
    .io_in_b(FP_multiplier_10ccs_31_io_in_b),
    .io_out_s(FP_multiplier_10ccs_31_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_32 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_32_clock),
    .reset(FP_multiplier_10ccs_32_reset),
    .io_in_a(FP_multiplier_10ccs_32_io_in_a),
    .io_in_b(FP_multiplier_10ccs_32_io_in_b),
    .io_out_s(FP_multiplier_10ccs_32_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_33 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_33_clock),
    .reset(FP_multiplier_10ccs_33_reset),
    .io_in_a(FP_multiplier_10ccs_33_io_in_a),
    .io_in_b(FP_multiplier_10ccs_33_io_in_b),
    .io_out_s(FP_multiplier_10ccs_33_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_34 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_34_clock),
    .reset(FP_multiplier_10ccs_34_reset),
    .io_in_a(FP_multiplier_10ccs_34_io_in_a),
    .io_in_b(FP_multiplier_10ccs_34_io_in_b),
    .io_out_s(FP_multiplier_10ccs_34_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_35 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_35_clock),
    .reset(FP_multiplier_10ccs_35_reset),
    .io_in_a(FP_multiplier_10ccs_35_io_in_a),
    .io_in_b(FP_multiplier_10ccs_35_io_in_b),
    .io_out_s(FP_multiplier_10ccs_35_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_36 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_36_clock),
    .reset(FP_multiplier_10ccs_36_reset),
    .io_in_a(FP_multiplier_10ccs_36_io_in_a),
    .io_in_b(FP_multiplier_10ccs_36_io_in_b),
    .io_out_s(FP_multiplier_10ccs_36_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_37 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_37_clock),
    .reset(FP_multiplier_10ccs_37_reset),
    .io_in_a(FP_multiplier_10ccs_37_io_in_a),
    .io_in_b(FP_multiplier_10ccs_37_io_in_b),
    .io_out_s(FP_multiplier_10ccs_37_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_38 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_38_clock),
    .reset(FP_multiplier_10ccs_38_reset),
    .io_in_a(FP_multiplier_10ccs_38_io_in_a),
    .io_in_b(FP_multiplier_10ccs_38_io_in_b),
    .io_out_s(FP_multiplier_10ccs_38_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_39 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_39_clock),
    .reset(FP_multiplier_10ccs_39_reset),
    .io_in_a(FP_multiplier_10ccs_39_io_in_a),
    .io_in_b(FP_multiplier_10ccs_39_io_in_b),
    .io_out_s(FP_multiplier_10ccs_39_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_40 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_40_clock),
    .reset(FP_multiplier_10ccs_40_reset),
    .io_in_a(FP_multiplier_10ccs_40_io_in_a),
    .io_in_b(FP_multiplier_10ccs_40_io_in_b),
    .io_out_s(FP_multiplier_10ccs_40_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_41 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_41_clock),
    .reset(FP_multiplier_10ccs_41_reset),
    .io_in_a(FP_multiplier_10ccs_41_io_in_a),
    .io_in_b(FP_multiplier_10ccs_41_io_in_b),
    .io_out_s(FP_multiplier_10ccs_41_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_42 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_42_clock),
    .reset(FP_multiplier_10ccs_42_reset),
    .io_in_a(FP_multiplier_10ccs_42_io_in_a),
    .io_in_b(FP_multiplier_10ccs_42_io_in_b),
    .io_out_s(FP_multiplier_10ccs_42_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_43 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_43_clock),
    .reset(FP_multiplier_10ccs_43_reset),
    .io_in_a(FP_multiplier_10ccs_43_io_in_a),
    .io_in_b(FP_multiplier_10ccs_43_io_in_b),
    .io_out_s(FP_multiplier_10ccs_43_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_44 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_44_clock),
    .reset(FP_multiplier_10ccs_44_reset),
    .io_in_a(FP_multiplier_10ccs_44_io_in_a),
    .io_in_b(FP_multiplier_10ccs_44_io_in_b),
    .io_out_s(FP_multiplier_10ccs_44_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_45 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_45_clock),
    .reset(FP_multiplier_10ccs_45_reset),
    .io_in_a(FP_multiplier_10ccs_45_io_in_a),
    .io_in_b(FP_multiplier_10ccs_45_io_in_b),
    .io_out_s(FP_multiplier_10ccs_45_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_46 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_46_clock),
    .reset(FP_multiplier_10ccs_46_reset),
    .io_in_a(FP_multiplier_10ccs_46_io_in_a),
    .io_in_b(FP_multiplier_10ccs_46_io_in_b),
    .io_out_s(FP_multiplier_10ccs_46_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_47 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_47_clock),
    .reset(FP_multiplier_10ccs_47_reset),
    .io_in_a(FP_multiplier_10ccs_47_io_in_a),
    .io_in_b(FP_multiplier_10ccs_47_io_in_b),
    .io_out_s(FP_multiplier_10ccs_47_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_48 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_48_clock),
    .reset(FP_multiplier_10ccs_48_reset),
    .io_in_a(FP_multiplier_10ccs_48_io_in_a),
    .io_in_b(FP_multiplier_10ccs_48_io_in_b),
    .io_out_s(FP_multiplier_10ccs_48_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_49 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_49_clock),
    .reset(FP_multiplier_10ccs_49_reset),
    .io_in_a(FP_multiplier_10ccs_49_io_in_a),
    .io_in_b(FP_multiplier_10ccs_49_io_in_b),
    .io_out_s(FP_multiplier_10ccs_49_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_50 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_50_clock),
    .reset(FP_multiplier_10ccs_50_reset),
    .io_in_a(FP_multiplier_10ccs_50_io_in_a),
    .io_in_b(FP_multiplier_10ccs_50_io_in_b),
    .io_out_s(FP_multiplier_10ccs_50_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_51 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_51_clock),
    .reset(FP_multiplier_10ccs_51_reset),
    .io_in_a(FP_multiplier_10ccs_51_io_in_a),
    .io_in_b(FP_multiplier_10ccs_51_io_in_b),
    .io_out_s(FP_multiplier_10ccs_51_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_52 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_52_clock),
    .reset(FP_multiplier_10ccs_52_reset),
    .io_in_a(FP_multiplier_10ccs_52_io_in_a),
    .io_in_b(FP_multiplier_10ccs_52_io_in_b),
    .io_out_s(FP_multiplier_10ccs_52_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_53 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_53_clock),
    .reset(FP_multiplier_10ccs_53_reset),
    .io_in_a(FP_multiplier_10ccs_53_io_in_a),
    .io_in_b(FP_multiplier_10ccs_53_io_in_b),
    .io_out_s(FP_multiplier_10ccs_53_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_54 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_54_clock),
    .reset(FP_multiplier_10ccs_54_reset),
    .io_in_a(FP_multiplier_10ccs_54_io_in_a),
    .io_in_b(FP_multiplier_10ccs_54_io_in_b),
    .io_out_s(FP_multiplier_10ccs_54_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_55 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_55_clock),
    .reset(FP_multiplier_10ccs_55_reset),
    .io_in_a(FP_multiplier_10ccs_55_io_in_a),
    .io_in_b(FP_multiplier_10ccs_55_io_in_b),
    .io_out_s(FP_multiplier_10ccs_55_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_56 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_56_clock),
    .reset(FP_multiplier_10ccs_56_reset),
    .io_in_a(FP_multiplier_10ccs_56_io_in_a),
    .io_in_b(FP_multiplier_10ccs_56_io_in_b),
    .io_out_s(FP_multiplier_10ccs_56_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_57 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_57_clock),
    .reset(FP_multiplier_10ccs_57_reset),
    .io_in_a(FP_multiplier_10ccs_57_io_in_a),
    .io_in_b(FP_multiplier_10ccs_57_io_in_b),
    .io_out_s(FP_multiplier_10ccs_57_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_58 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_58_clock),
    .reset(FP_multiplier_10ccs_58_reset),
    .io_in_a(FP_multiplier_10ccs_58_io_in_a),
    .io_in_b(FP_multiplier_10ccs_58_io_in_b),
    .io_out_s(FP_multiplier_10ccs_58_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_59 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_59_clock),
    .reset(FP_multiplier_10ccs_59_reset),
    .io_in_a(FP_multiplier_10ccs_59_io_in_a),
    .io_in_b(FP_multiplier_10ccs_59_io_in_b),
    .io_out_s(FP_multiplier_10ccs_59_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_60 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_60_clock),
    .reset(FP_multiplier_10ccs_60_reset),
    .io_in_a(FP_multiplier_10ccs_60_io_in_a),
    .io_in_b(FP_multiplier_10ccs_60_io_in_b),
    .io_out_s(FP_multiplier_10ccs_60_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_61 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_61_clock),
    .reset(FP_multiplier_10ccs_61_reset),
    .io_in_a(FP_multiplier_10ccs_61_io_in_a),
    .io_in_b(FP_multiplier_10ccs_61_io_in_b),
    .io_out_s(FP_multiplier_10ccs_61_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_62 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_62_clock),
    .reset(FP_multiplier_10ccs_62_reset),
    .io_in_a(FP_multiplier_10ccs_62_io_in_a),
    .io_in_b(FP_multiplier_10ccs_62_io_in_b),
    .io_out_s(FP_multiplier_10ccs_62_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_63 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_63_clock),
    .reset(FP_multiplier_10ccs_63_reset),
    .io_in_a(FP_multiplier_10ccs_63_io_in_a),
    .io_in_b(FP_multiplier_10ccs_63_io_in_b),
    .io_out_s(FP_multiplier_10ccs_63_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_64 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_64_clock),
    .reset(FP_multiplier_10ccs_64_reset),
    .io_in_a(FP_multiplier_10ccs_64_io_in_a),
    .io_in_b(FP_multiplier_10ccs_64_io_in_b),
    .io_out_s(FP_multiplier_10ccs_64_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_65 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_65_clock),
    .reset(FP_multiplier_10ccs_65_reset),
    .io_in_a(FP_multiplier_10ccs_65_io_in_a),
    .io_in_b(FP_multiplier_10ccs_65_io_in_b),
    .io_out_s(FP_multiplier_10ccs_65_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_66 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_66_clock),
    .reset(FP_multiplier_10ccs_66_reset),
    .io_in_a(FP_multiplier_10ccs_66_io_in_a),
    .io_in_b(FP_multiplier_10ccs_66_io_in_b),
    .io_out_s(FP_multiplier_10ccs_66_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_67 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_67_clock),
    .reset(FP_multiplier_10ccs_67_reset),
    .io_in_a(FP_multiplier_10ccs_67_io_in_a),
    .io_in_b(FP_multiplier_10ccs_67_io_in_b),
    .io_out_s(FP_multiplier_10ccs_67_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_68 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_68_clock),
    .reset(FP_multiplier_10ccs_68_reset),
    .io_in_a(FP_multiplier_10ccs_68_io_in_a),
    .io_in_b(FP_multiplier_10ccs_68_io_in_b),
    .io_out_s(FP_multiplier_10ccs_68_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_69 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_69_clock),
    .reset(FP_multiplier_10ccs_69_reset),
    .io_in_a(FP_multiplier_10ccs_69_io_in_a),
    .io_in_b(FP_multiplier_10ccs_69_io_in_b),
    .io_out_s(FP_multiplier_10ccs_69_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_70 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_70_clock),
    .reset(FP_multiplier_10ccs_70_reset),
    .io_in_a(FP_multiplier_10ccs_70_io_in_a),
    .io_in_b(FP_multiplier_10ccs_70_io_in_b),
    .io_out_s(FP_multiplier_10ccs_70_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_71 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_71_clock),
    .reset(FP_multiplier_10ccs_71_reset),
    .io_in_a(FP_multiplier_10ccs_71_io_in_a),
    .io_in_b(FP_multiplier_10ccs_71_io_in_b),
    .io_out_s(FP_multiplier_10ccs_71_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_72 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_72_clock),
    .reset(FP_multiplier_10ccs_72_reset),
    .io_in_a(FP_multiplier_10ccs_72_io_in_a),
    .io_in_b(FP_multiplier_10ccs_72_io_in_b),
    .io_out_s(FP_multiplier_10ccs_72_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_73 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_73_clock),
    .reset(FP_multiplier_10ccs_73_reset),
    .io_in_a(FP_multiplier_10ccs_73_io_in_a),
    .io_in_b(FP_multiplier_10ccs_73_io_in_b),
    .io_out_s(FP_multiplier_10ccs_73_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_74 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_74_clock),
    .reset(FP_multiplier_10ccs_74_reset),
    .io_in_a(FP_multiplier_10ccs_74_io_in_a),
    .io_in_b(FP_multiplier_10ccs_74_io_in_b),
    .io_out_s(FP_multiplier_10ccs_74_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_75 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_75_clock),
    .reset(FP_multiplier_10ccs_75_reset),
    .io_in_a(FP_multiplier_10ccs_75_io_in_a),
    .io_in_b(FP_multiplier_10ccs_75_io_in_b),
    .io_out_s(FP_multiplier_10ccs_75_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_76 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_76_clock),
    .reset(FP_multiplier_10ccs_76_reset),
    .io_in_a(FP_multiplier_10ccs_76_io_in_a),
    .io_in_b(FP_multiplier_10ccs_76_io_in_b),
    .io_out_s(FP_multiplier_10ccs_76_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_77 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_77_clock),
    .reset(FP_multiplier_10ccs_77_reset),
    .io_in_a(FP_multiplier_10ccs_77_io_in_a),
    .io_in_b(FP_multiplier_10ccs_77_io_in_b),
    .io_out_s(FP_multiplier_10ccs_77_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_78 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_78_clock),
    .reset(FP_multiplier_10ccs_78_reset),
    .io_in_a(FP_multiplier_10ccs_78_io_in_a),
    .io_in_b(FP_multiplier_10ccs_78_io_in_b),
    .io_out_s(FP_multiplier_10ccs_78_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_79 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_79_clock),
    .reset(FP_multiplier_10ccs_79_reset),
    .io_in_a(FP_multiplier_10ccs_79_io_in_a),
    .io_in_b(FP_multiplier_10ccs_79_io_in_b),
    .io_out_s(FP_multiplier_10ccs_79_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_80 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_80_clock),
    .reset(FP_multiplier_10ccs_80_reset),
    .io_in_a(FP_multiplier_10ccs_80_io_in_a),
    .io_in_b(FP_multiplier_10ccs_80_io_in_b),
    .io_out_s(FP_multiplier_10ccs_80_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_81 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_81_clock),
    .reset(FP_multiplier_10ccs_81_reset),
    .io_in_a(FP_multiplier_10ccs_81_io_in_a),
    .io_in_b(FP_multiplier_10ccs_81_io_in_b),
    .io_out_s(FP_multiplier_10ccs_81_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_82 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_82_clock),
    .reset(FP_multiplier_10ccs_82_reset),
    .io_in_a(FP_multiplier_10ccs_82_io_in_a),
    .io_in_b(FP_multiplier_10ccs_82_io_in_b),
    .io_out_s(FP_multiplier_10ccs_82_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_83 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_83_clock),
    .reset(FP_multiplier_10ccs_83_reset),
    .io_in_a(FP_multiplier_10ccs_83_io_in_a),
    .io_in_b(FP_multiplier_10ccs_83_io_in_b),
    .io_out_s(FP_multiplier_10ccs_83_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_84 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_84_clock),
    .reset(FP_multiplier_10ccs_84_reset),
    .io_in_a(FP_multiplier_10ccs_84_io_in_a),
    .io_in_b(FP_multiplier_10ccs_84_io_in_b),
    .io_out_s(FP_multiplier_10ccs_84_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_85 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_85_clock),
    .reset(FP_multiplier_10ccs_85_reset),
    .io_in_a(FP_multiplier_10ccs_85_io_in_a),
    .io_in_b(FP_multiplier_10ccs_85_io_in_b),
    .io_out_s(FP_multiplier_10ccs_85_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_86 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_86_clock),
    .reset(FP_multiplier_10ccs_86_reset),
    .io_in_a(FP_multiplier_10ccs_86_io_in_a),
    .io_in_b(FP_multiplier_10ccs_86_io_in_b),
    .io_out_s(FP_multiplier_10ccs_86_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_87 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_87_clock),
    .reset(FP_multiplier_10ccs_87_reset),
    .io_in_a(FP_multiplier_10ccs_87_io_in_a),
    .io_in_b(FP_multiplier_10ccs_87_io_in_b),
    .io_out_s(FP_multiplier_10ccs_87_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_88 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_88_clock),
    .reset(FP_multiplier_10ccs_88_reset),
    .io_in_a(FP_multiplier_10ccs_88_io_in_a),
    .io_in_b(FP_multiplier_10ccs_88_io_in_b),
    .io_out_s(FP_multiplier_10ccs_88_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_89 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_89_clock),
    .reset(FP_multiplier_10ccs_89_reset),
    .io_in_a(FP_multiplier_10ccs_89_io_in_a),
    .io_in_b(FP_multiplier_10ccs_89_io_in_b),
    .io_out_s(FP_multiplier_10ccs_89_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_90 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_90_clock),
    .reset(FP_multiplier_10ccs_90_reset),
    .io_in_a(FP_multiplier_10ccs_90_io_in_a),
    .io_in_b(FP_multiplier_10ccs_90_io_in_b),
    .io_out_s(FP_multiplier_10ccs_90_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_91 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_91_clock),
    .reset(FP_multiplier_10ccs_91_reset),
    .io_in_a(FP_multiplier_10ccs_91_io_in_a),
    .io_in_b(FP_multiplier_10ccs_91_io_in_b),
    .io_out_s(FP_multiplier_10ccs_91_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_92 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_92_clock),
    .reset(FP_multiplier_10ccs_92_reset),
    .io_in_a(FP_multiplier_10ccs_92_io_in_a),
    .io_in_b(FP_multiplier_10ccs_92_io_in_b),
    .io_out_s(FP_multiplier_10ccs_92_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_93 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_93_clock),
    .reset(FP_multiplier_10ccs_93_reset),
    .io_in_a(FP_multiplier_10ccs_93_io_in_a),
    .io_in_b(FP_multiplier_10ccs_93_io_in_b),
    .io_out_s(FP_multiplier_10ccs_93_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_94 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_94_clock),
    .reset(FP_multiplier_10ccs_94_reset),
    .io_in_a(FP_multiplier_10ccs_94_io_in_a),
    .io_in_b(FP_multiplier_10ccs_94_io_in_b),
    .io_out_s(FP_multiplier_10ccs_94_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_95 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_95_clock),
    .reset(FP_multiplier_10ccs_95_reset),
    .io_in_a(FP_multiplier_10ccs_95_io_in_a),
    .io_in_b(FP_multiplier_10ccs_95_io_in_b),
    .io_out_s(FP_multiplier_10ccs_95_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_96 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_96_clock),
    .reset(FP_multiplier_10ccs_96_reset),
    .io_in_a(FP_multiplier_10ccs_96_io_in_a),
    .io_in_b(FP_multiplier_10ccs_96_io_in_b),
    .io_out_s(FP_multiplier_10ccs_96_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_97 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_97_clock),
    .reset(FP_multiplier_10ccs_97_reset),
    .io_in_a(FP_multiplier_10ccs_97_io_in_a),
    .io_in_b(FP_multiplier_10ccs_97_io_in_b),
    .io_out_s(FP_multiplier_10ccs_97_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_98 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_98_clock),
    .reset(FP_multiplier_10ccs_98_reset),
    .io_in_a(FP_multiplier_10ccs_98_io_in_a),
    .io_in_b(FP_multiplier_10ccs_98_io_in_b),
    .io_out_s(FP_multiplier_10ccs_98_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_99 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_99_clock),
    .reset(FP_multiplier_10ccs_99_reset),
    .io_in_a(FP_multiplier_10ccs_99_io_in_a),
    .io_in_b(FP_multiplier_10ccs_99_io_in_b),
    .io_out_s(FP_multiplier_10ccs_99_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_100 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_100_clock),
    .reset(FP_multiplier_10ccs_100_reset),
    .io_in_a(FP_multiplier_10ccs_100_io_in_a),
    .io_in_b(FP_multiplier_10ccs_100_io_in_b),
    .io_out_s(FP_multiplier_10ccs_100_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_101 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_101_clock),
    .reset(FP_multiplier_10ccs_101_reset),
    .io_in_a(FP_multiplier_10ccs_101_io_in_a),
    .io_in_b(FP_multiplier_10ccs_101_io_in_b),
    .io_out_s(FP_multiplier_10ccs_101_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_102 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_102_clock),
    .reset(FP_multiplier_10ccs_102_reset),
    .io_in_a(FP_multiplier_10ccs_102_io_in_a),
    .io_in_b(FP_multiplier_10ccs_102_io_in_b),
    .io_out_s(FP_multiplier_10ccs_102_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_103 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_103_clock),
    .reset(FP_multiplier_10ccs_103_reset),
    .io_in_a(FP_multiplier_10ccs_103_io_in_a),
    .io_in_b(FP_multiplier_10ccs_103_io_in_b),
    .io_out_s(FP_multiplier_10ccs_103_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_104 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_104_clock),
    .reset(FP_multiplier_10ccs_104_reset),
    .io_in_a(FP_multiplier_10ccs_104_io_in_a),
    .io_in_b(FP_multiplier_10ccs_104_io_in_b),
    .io_out_s(FP_multiplier_10ccs_104_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_105 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_105_clock),
    .reset(FP_multiplier_10ccs_105_reset),
    .io_in_a(FP_multiplier_10ccs_105_io_in_a),
    .io_in_b(FP_multiplier_10ccs_105_io_in_b),
    .io_out_s(FP_multiplier_10ccs_105_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_106 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_106_clock),
    .reset(FP_multiplier_10ccs_106_reset),
    .io_in_a(FP_multiplier_10ccs_106_io_in_a),
    .io_in_b(FP_multiplier_10ccs_106_io_in_b),
    .io_out_s(FP_multiplier_10ccs_106_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_107 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_107_clock),
    .reset(FP_multiplier_10ccs_107_reset),
    .io_in_a(FP_multiplier_10ccs_107_io_in_a),
    .io_in_b(FP_multiplier_10ccs_107_io_in_b),
    .io_out_s(FP_multiplier_10ccs_107_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_108 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_108_clock),
    .reset(FP_multiplier_10ccs_108_reset),
    .io_in_a(FP_multiplier_10ccs_108_io_in_a),
    .io_in_b(FP_multiplier_10ccs_108_io_in_b),
    .io_out_s(FP_multiplier_10ccs_108_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_109 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_109_clock),
    .reset(FP_multiplier_10ccs_109_reset),
    .io_in_a(FP_multiplier_10ccs_109_io_in_a),
    .io_in_b(FP_multiplier_10ccs_109_io_in_b),
    .io_out_s(FP_multiplier_10ccs_109_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_110 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_110_clock),
    .reset(FP_multiplier_10ccs_110_reset),
    .io_in_a(FP_multiplier_10ccs_110_io_in_a),
    .io_in_b(FP_multiplier_10ccs_110_io_in_b),
    .io_out_s(FP_multiplier_10ccs_110_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_111 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_111_clock),
    .reset(FP_multiplier_10ccs_111_reset),
    .io_in_a(FP_multiplier_10ccs_111_io_in_a),
    .io_in_b(FP_multiplier_10ccs_111_io_in_b),
    .io_out_s(FP_multiplier_10ccs_111_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_112 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_112_clock),
    .reset(FP_multiplier_10ccs_112_reset),
    .io_in_a(FP_multiplier_10ccs_112_io_in_a),
    .io_in_b(FP_multiplier_10ccs_112_io_in_b),
    .io_out_s(FP_multiplier_10ccs_112_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_113 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_113_clock),
    .reset(FP_multiplier_10ccs_113_reset),
    .io_in_a(FP_multiplier_10ccs_113_io_in_a),
    .io_in_b(FP_multiplier_10ccs_113_io_in_b),
    .io_out_s(FP_multiplier_10ccs_113_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_114 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_114_clock),
    .reset(FP_multiplier_10ccs_114_reset),
    .io_in_a(FP_multiplier_10ccs_114_io_in_a),
    .io_in_b(FP_multiplier_10ccs_114_io_in_b),
    .io_out_s(FP_multiplier_10ccs_114_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_115 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_115_clock),
    .reset(FP_multiplier_10ccs_115_reset),
    .io_in_a(FP_multiplier_10ccs_115_io_in_a),
    .io_in_b(FP_multiplier_10ccs_115_io_in_b),
    .io_out_s(FP_multiplier_10ccs_115_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_116 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_116_clock),
    .reset(FP_multiplier_10ccs_116_reset),
    .io_in_a(FP_multiplier_10ccs_116_io_in_a),
    .io_in_b(FP_multiplier_10ccs_116_io_in_b),
    .io_out_s(FP_multiplier_10ccs_116_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_117 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_117_clock),
    .reset(FP_multiplier_10ccs_117_reset),
    .io_in_a(FP_multiplier_10ccs_117_io_in_a),
    .io_in_b(FP_multiplier_10ccs_117_io_in_b),
    .io_out_s(FP_multiplier_10ccs_117_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_118 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_118_clock),
    .reset(FP_multiplier_10ccs_118_reset),
    .io_in_a(FP_multiplier_10ccs_118_io_in_a),
    .io_in_b(FP_multiplier_10ccs_118_io_in_b),
    .io_out_s(FP_multiplier_10ccs_118_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_119 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_119_clock),
    .reset(FP_multiplier_10ccs_119_reset),
    .io_in_a(FP_multiplier_10ccs_119_io_in_a),
    .io_in_b(FP_multiplier_10ccs_119_io_in_b),
    .io_out_s(FP_multiplier_10ccs_119_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_120 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_120_clock),
    .reset(FP_multiplier_10ccs_120_reset),
    .io_in_a(FP_multiplier_10ccs_120_io_in_a),
    .io_in_b(FP_multiplier_10ccs_120_io_in_b),
    .io_out_s(FP_multiplier_10ccs_120_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_121 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_121_clock),
    .reset(FP_multiplier_10ccs_121_reset),
    .io_in_a(FP_multiplier_10ccs_121_io_in_a),
    .io_in_b(FP_multiplier_10ccs_121_io_in_b),
    .io_out_s(FP_multiplier_10ccs_121_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_122 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_122_clock),
    .reset(FP_multiplier_10ccs_122_reset),
    .io_in_a(FP_multiplier_10ccs_122_io_in_a),
    .io_in_b(FP_multiplier_10ccs_122_io_in_b),
    .io_out_s(FP_multiplier_10ccs_122_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_123 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_123_clock),
    .reset(FP_multiplier_10ccs_123_reset),
    .io_in_a(FP_multiplier_10ccs_123_io_in_a),
    .io_in_b(FP_multiplier_10ccs_123_io_in_b),
    .io_out_s(FP_multiplier_10ccs_123_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_124 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_124_clock),
    .reset(FP_multiplier_10ccs_124_reset),
    .io_in_a(FP_multiplier_10ccs_124_io_in_a),
    .io_in_b(FP_multiplier_10ccs_124_io_in_b),
    .io_out_s(FP_multiplier_10ccs_124_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_125 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_125_clock),
    .reset(FP_multiplier_10ccs_125_reset),
    .io_in_a(FP_multiplier_10ccs_125_io_in_a),
    .io_in_b(FP_multiplier_10ccs_125_io_in_b),
    .io_out_s(FP_multiplier_10ccs_125_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_126 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_126_clock),
    .reset(FP_multiplier_10ccs_126_reset),
    .io_in_a(FP_multiplier_10ccs_126_io_in_a),
    .io_in_b(FP_multiplier_10ccs_126_io_in_b),
    .io_out_s(FP_multiplier_10ccs_126_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_127 ( // @[FloatingPointDesigns.scala 2483:28]
    .clock(FP_multiplier_10ccs_127_clock),
    .reset(FP_multiplier_10ccs_127_reset),
    .io_in_a(FP_multiplier_10ccs_127_io_in_a),
    .io_in_b(FP_multiplier_10ccs_127_io_in_b),
    .io_out_s(FP_multiplier_10ccs_127_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_clock),
    .reset(FP_adder_13ccs_reset),
    .io_in_a(FP_adder_13ccs_io_in_a),
    .io_in_b(FP_adder_13ccs_io_in_b),
    .io_out_s(FP_adder_13ccs_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_1 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_1_clock),
    .reset(FP_adder_13ccs_1_reset),
    .io_in_a(FP_adder_13ccs_1_io_in_a),
    .io_in_b(FP_adder_13ccs_1_io_in_b),
    .io_out_s(FP_adder_13ccs_1_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_2 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_2_clock),
    .reset(FP_adder_13ccs_2_reset),
    .io_in_a(FP_adder_13ccs_2_io_in_a),
    .io_in_b(FP_adder_13ccs_2_io_in_b),
    .io_out_s(FP_adder_13ccs_2_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_3 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_3_clock),
    .reset(FP_adder_13ccs_3_reset),
    .io_in_a(FP_adder_13ccs_3_io_in_a),
    .io_in_b(FP_adder_13ccs_3_io_in_b),
    .io_out_s(FP_adder_13ccs_3_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_4 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_4_clock),
    .reset(FP_adder_13ccs_4_reset),
    .io_in_a(FP_adder_13ccs_4_io_in_a),
    .io_in_b(FP_adder_13ccs_4_io_in_b),
    .io_out_s(FP_adder_13ccs_4_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_5 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_5_clock),
    .reset(FP_adder_13ccs_5_reset),
    .io_in_a(FP_adder_13ccs_5_io_in_a),
    .io_in_b(FP_adder_13ccs_5_io_in_b),
    .io_out_s(FP_adder_13ccs_5_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_6 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_6_clock),
    .reset(FP_adder_13ccs_6_reset),
    .io_in_a(FP_adder_13ccs_6_io_in_a),
    .io_in_b(FP_adder_13ccs_6_io_in_b),
    .io_out_s(FP_adder_13ccs_6_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_7 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_7_clock),
    .reset(FP_adder_13ccs_7_reset),
    .io_in_a(FP_adder_13ccs_7_io_in_a),
    .io_in_b(FP_adder_13ccs_7_io_in_b),
    .io_out_s(FP_adder_13ccs_7_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_8 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_8_clock),
    .reset(FP_adder_13ccs_8_reset),
    .io_in_a(FP_adder_13ccs_8_io_in_a),
    .io_in_b(FP_adder_13ccs_8_io_in_b),
    .io_out_s(FP_adder_13ccs_8_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_9 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_9_clock),
    .reset(FP_adder_13ccs_9_reset),
    .io_in_a(FP_adder_13ccs_9_io_in_a),
    .io_in_b(FP_adder_13ccs_9_io_in_b),
    .io_out_s(FP_adder_13ccs_9_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_10 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_10_clock),
    .reset(FP_adder_13ccs_10_reset),
    .io_in_a(FP_adder_13ccs_10_io_in_a),
    .io_in_b(FP_adder_13ccs_10_io_in_b),
    .io_out_s(FP_adder_13ccs_10_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_11 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_11_clock),
    .reset(FP_adder_13ccs_11_reset),
    .io_in_a(FP_adder_13ccs_11_io_in_a),
    .io_in_b(FP_adder_13ccs_11_io_in_b),
    .io_out_s(FP_adder_13ccs_11_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_12 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_12_clock),
    .reset(FP_adder_13ccs_12_reset),
    .io_in_a(FP_adder_13ccs_12_io_in_a),
    .io_in_b(FP_adder_13ccs_12_io_in_b),
    .io_out_s(FP_adder_13ccs_12_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_13 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_13_clock),
    .reset(FP_adder_13ccs_13_reset),
    .io_in_a(FP_adder_13ccs_13_io_in_a),
    .io_in_b(FP_adder_13ccs_13_io_in_b),
    .io_out_s(FP_adder_13ccs_13_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_14 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_14_clock),
    .reset(FP_adder_13ccs_14_reset),
    .io_in_a(FP_adder_13ccs_14_io_in_a),
    .io_in_b(FP_adder_13ccs_14_io_in_b),
    .io_out_s(FP_adder_13ccs_14_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_15 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_15_clock),
    .reset(FP_adder_13ccs_15_reset),
    .io_in_a(FP_adder_13ccs_15_io_in_a),
    .io_in_b(FP_adder_13ccs_15_io_in_b),
    .io_out_s(FP_adder_13ccs_15_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_16 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_16_clock),
    .reset(FP_adder_13ccs_16_reset),
    .io_in_a(FP_adder_13ccs_16_io_in_a),
    .io_in_b(FP_adder_13ccs_16_io_in_b),
    .io_out_s(FP_adder_13ccs_16_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_17 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_17_clock),
    .reset(FP_adder_13ccs_17_reset),
    .io_in_a(FP_adder_13ccs_17_io_in_a),
    .io_in_b(FP_adder_13ccs_17_io_in_b),
    .io_out_s(FP_adder_13ccs_17_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_18 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_18_clock),
    .reset(FP_adder_13ccs_18_reset),
    .io_in_a(FP_adder_13ccs_18_io_in_a),
    .io_in_b(FP_adder_13ccs_18_io_in_b),
    .io_out_s(FP_adder_13ccs_18_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_19 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_19_clock),
    .reset(FP_adder_13ccs_19_reset),
    .io_in_a(FP_adder_13ccs_19_io_in_a),
    .io_in_b(FP_adder_13ccs_19_io_in_b),
    .io_out_s(FP_adder_13ccs_19_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_20 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_20_clock),
    .reset(FP_adder_13ccs_20_reset),
    .io_in_a(FP_adder_13ccs_20_io_in_a),
    .io_in_b(FP_adder_13ccs_20_io_in_b),
    .io_out_s(FP_adder_13ccs_20_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_21 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_21_clock),
    .reset(FP_adder_13ccs_21_reset),
    .io_in_a(FP_adder_13ccs_21_io_in_a),
    .io_in_b(FP_adder_13ccs_21_io_in_b),
    .io_out_s(FP_adder_13ccs_21_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_22 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_22_clock),
    .reset(FP_adder_13ccs_22_reset),
    .io_in_a(FP_adder_13ccs_22_io_in_a),
    .io_in_b(FP_adder_13ccs_22_io_in_b),
    .io_out_s(FP_adder_13ccs_22_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_23 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_23_clock),
    .reset(FP_adder_13ccs_23_reset),
    .io_in_a(FP_adder_13ccs_23_io_in_a),
    .io_in_b(FP_adder_13ccs_23_io_in_b),
    .io_out_s(FP_adder_13ccs_23_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_24 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_24_clock),
    .reset(FP_adder_13ccs_24_reset),
    .io_in_a(FP_adder_13ccs_24_io_in_a),
    .io_in_b(FP_adder_13ccs_24_io_in_b),
    .io_out_s(FP_adder_13ccs_24_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_25 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_25_clock),
    .reset(FP_adder_13ccs_25_reset),
    .io_in_a(FP_adder_13ccs_25_io_in_a),
    .io_in_b(FP_adder_13ccs_25_io_in_b),
    .io_out_s(FP_adder_13ccs_25_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_26 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_26_clock),
    .reset(FP_adder_13ccs_26_reset),
    .io_in_a(FP_adder_13ccs_26_io_in_a),
    .io_in_b(FP_adder_13ccs_26_io_in_b),
    .io_out_s(FP_adder_13ccs_26_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_27 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_27_clock),
    .reset(FP_adder_13ccs_27_reset),
    .io_in_a(FP_adder_13ccs_27_io_in_a),
    .io_in_b(FP_adder_13ccs_27_io_in_b),
    .io_out_s(FP_adder_13ccs_27_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_28 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_28_clock),
    .reset(FP_adder_13ccs_28_reset),
    .io_in_a(FP_adder_13ccs_28_io_in_a),
    .io_in_b(FP_adder_13ccs_28_io_in_b),
    .io_out_s(FP_adder_13ccs_28_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_29 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_29_clock),
    .reset(FP_adder_13ccs_29_reset),
    .io_in_a(FP_adder_13ccs_29_io_in_a),
    .io_in_b(FP_adder_13ccs_29_io_in_b),
    .io_out_s(FP_adder_13ccs_29_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_30 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_30_clock),
    .reset(FP_adder_13ccs_30_reset),
    .io_in_a(FP_adder_13ccs_30_io_in_a),
    .io_in_b(FP_adder_13ccs_30_io_in_b),
    .io_out_s(FP_adder_13ccs_30_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_31 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_31_clock),
    .reset(FP_adder_13ccs_31_reset),
    .io_in_a(FP_adder_13ccs_31_io_in_a),
    .io_in_b(FP_adder_13ccs_31_io_in_b),
    .io_out_s(FP_adder_13ccs_31_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_32 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_32_clock),
    .reset(FP_adder_13ccs_32_reset),
    .io_in_a(FP_adder_13ccs_32_io_in_a),
    .io_in_b(FP_adder_13ccs_32_io_in_b),
    .io_out_s(FP_adder_13ccs_32_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_33 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_33_clock),
    .reset(FP_adder_13ccs_33_reset),
    .io_in_a(FP_adder_13ccs_33_io_in_a),
    .io_in_b(FP_adder_13ccs_33_io_in_b),
    .io_out_s(FP_adder_13ccs_33_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_34 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_34_clock),
    .reset(FP_adder_13ccs_34_reset),
    .io_in_a(FP_adder_13ccs_34_io_in_a),
    .io_in_b(FP_adder_13ccs_34_io_in_b),
    .io_out_s(FP_adder_13ccs_34_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_35 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_35_clock),
    .reset(FP_adder_13ccs_35_reset),
    .io_in_a(FP_adder_13ccs_35_io_in_a),
    .io_in_b(FP_adder_13ccs_35_io_in_b),
    .io_out_s(FP_adder_13ccs_35_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_36 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_36_clock),
    .reset(FP_adder_13ccs_36_reset),
    .io_in_a(FP_adder_13ccs_36_io_in_a),
    .io_in_b(FP_adder_13ccs_36_io_in_b),
    .io_out_s(FP_adder_13ccs_36_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_37 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_37_clock),
    .reset(FP_adder_13ccs_37_reset),
    .io_in_a(FP_adder_13ccs_37_io_in_a),
    .io_in_b(FP_adder_13ccs_37_io_in_b),
    .io_out_s(FP_adder_13ccs_37_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_38 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_38_clock),
    .reset(FP_adder_13ccs_38_reset),
    .io_in_a(FP_adder_13ccs_38_io_in_a),
    .io_in_b(FP_adder_13ccs_38_io_in_b),
    .io_out_s(FP_adder_13ccs_38_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_39 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_39_clock),
    .reset(FP_adder_13ccs_39_reset),
    .io_in_a(FP_adder_13ccs_39_io_in_a),
    .io_in_b(FP_adder_13ccs_39_io_in_b),
    .io_out_s(FP_adder_13ccs_39_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_40 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_40_clock),
    .reset(FP_adder_13ccs_40_reset),
    .io_in_a(FP_adder_13ccs_40_io_in_a),
    .io_in_b(FP_adder_13ccs_40_io_in_b),
    .io_out_s(FP_adder_13ccs_40_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_41 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_41_clock),
    .reset(FP_adder_13ccs_41_reset),
    .io_in_a(FP_adder_13ccs_41_io_in_a),
    .io_in_b(FP_adder_13ccs_41_io_in_b),
    .io_out_s(FP_adder_13ccs_41_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_42 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_42_clock),
    .reset(FP_adder_13ccs_42_reset),
    .io_in_a(FP_adder_13ccs_42_io_in_a),
    .io_in_b(FP_adder_13ccs_42_io_in_b),
    .io_out_s(FP_adder_13ccs_42_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_43 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_43_clock),
    .reset(FP_adder_13ccs_43_reset),
    .io_in_a(FP_adder_13ccs_43_io_in_a),
    .io_in_b(FP_adder_13ccs_43_io_in_b),
    .io_out_s(FP_adder_13ccs_43_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_44 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_44_clock),
    .reset(FP_adder_13ccs_44_reset),
    .io_in_a(FP_adder_13ccs_44_io_in_a),
    .io_in_b(FP_adder_13ccs_44_io_in_b),
    .io_out_s(FP_adder_13ccs_44_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_45 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_45_clock),
    .reset(FP_adder_13ccs_45_reset),
    .io_in_a(FP_adder_13ccs_45_io_in_a),
    .io_in_b(FP_adder_13ccs_45_io_in_b),
    .io_out_s(FP_adder_13ccs_45_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_46 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_46_clock),
    .reset(FP_adder_13ccs_46_reset),
    .io_in_a(FP_adder_13ccs_46_io_in_a),
    .io_in_b(FP_adder_13ccs_46_io_in_b),
    .io_out_s(FP_adder_13ccs_46_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_47 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_47_clock),
    .reset(FP_adder_13ccs_47_reset),
    .io_in_a(FP_adder_13ccs_47_io_in_a),
    .io_in_b(FP_adder_13ccs_47_io_in_b),
    .io_out_s(FP_adder_13ccs_47_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_48 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_48_clock),
    .reset(FP_adder_13ccs_48_reset),
    .io_in_a(FP_adder_13ccs_48_io_in_a),
    .io_in_b(FP_adder_13ccs_48_io_in_b),
    .io_out_s(FP_adder_13ccs_48_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_49 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_49_clock),
    .reset(FP_adder_13ccs_49_reset),
    .io_in_a(FP_adder_13ccs_49_io_in_a),
    .io_in_b(FP_adder_13ccs_49_io_in_b),
    .io_out_s(FP_adder_13ccs_49_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_50 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_50_clock),
    .reset(FP_adder_13ccs_50_reset),
    .io_in_a(FP_adder_13ccs_50_io_in_a),
    .io_in_b(FP_adder_13ccs_50_io_in_b),
    .io_out_s(FP_adder_13ccs_50_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_51 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_51_clock),
    .reset(FP_adder_13ccs_51_reset),
    .io_in_a(FP_adder_13ccs_51_io_in_a),
    .io_in_b(FP_adder_13ccs_51_io_in_b),
    .io_out_s(FP_adder_13ccs_51_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_52 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_52_clock),
    .reset(FP_adder_13ccs_52_reset),
    .io_in_a(FP_adder_13ccs_52_io_in_a),
    .io_in_b(FP_adder_13ccs_52_io_in_b),
    .io_out_s(FP_adder_13ccs_52_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_53 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_53_clock),
    .reset(FP_adder_13ccs_53_reset),
    .io_in_a(FP_adder_13ccs_53_io_in_a),
    .io_in_b(FP_adder_13ccs_53_io_in_b),
    .io_out_s(FP_adder_13ccs_53_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_54 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_54_clock),
    .reset(FP_adder_13ccs_54_reset),
    .io_in_a(FP_adder_13ccs_54_io_in_a),
    .io_in_b(FP_adder_13ccs_54_io_in_b),
    .io_out_s(FP_adder_13ccs_54_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_55 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_55_clock),
    .reset(FP_adder_13ccs_55_reset),
    .io_in_a(FP_adder_13ccs_55_io_in_a),
    .io_in_b(FP_adder_13ccs_55_io_in_b),
    .io_out_s(FP_adder_13ccs_55_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_56 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_56_clock),
    .reset(FP_adder_13ccs_56_reset),
    .io_in_a(FP_adder_13ccs_56_io_in_a),
    .io_in_b(FP_adder_13ccs_56_io_in_b),
    .io_out_s(FP_adder_13ccs_56_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_57 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_57_clock),
    .reset(FP_adder_13ccs_57_reset),
    .io_in_a(FP_adder_13ccs_57_io_in_a),
    .io_in_b(FP_adder_13ccs_57_io_in_b),
    .io_out_s(FP_adder_13ccs_57_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_58 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_58_clock),
    .reset(FP_adder_13ccs_58_reset),
    .io_in_a(FP_adder_13ccs_58_io_in_a),
    .io_in_b(FP_adder_13ccs_58_io_in_b),
    .io_out_s(FP_adder_13ccs_58_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_59 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_59_clock),
    .reset(FP_adder_13ccs_59_reset),
    .io_in_a(FP_adder_13ccs_59_io_in_a),
    .io_in_b(FP_adder_13ccs_59_io_in_b),
    .io_out_s(FP_adder_13ccs_59_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_60 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_60_clock),
    .reset(FP_adder_13ccs_60_reset),
    .io_in_a(FP_adder_13ccs_60_io_in_a),
    .io_in_b(FP_adder_13ccs_60_io_in_b),
    .io_out_s(FP_adder_13ccs_60_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_61 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_61_clock),
    .reset(FP_adder_13ccs_61_reset),
    .io_in_a(FP_adder_13ccs_61_io_in_a),
    .io_in_b(FP_adder_13ccs_61_io_in_b),
    .io_out_s(FP_adder_13ccs_61_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_62 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_62_clock),
    .reset(FP_adder_13ccs_62_reset),
    .io_in_a(FP_adder_13ccs_62_io_in_a),
    .io_in_b(FP_adder_13ccs_62_io_in_b),
    .io_out_s(FP_adder_13ccs_62_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_63 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_63_clock),
    .reset(FP_adder_13ccs_63_reset),
    .io_in_a(FP_adder_13ccs_63_io_in_a),
    .io_in_b(FP_adder_13ccs_63_io_in_b),
    .io_out_s(FP_adder_13ccs_63_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_64 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_64_clock),
    .reset(FP_adder_13ccs_64_reset),
    .io_in_a(FP_adder_13ccs_64_io_in_a),
    .io_in_b(FP_adder_13ccs_64_io_in_b),
    .io_out_s(FP_adder_13ccs_64_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_65 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_65_clock),
    .reset(FP_adder_13ccs_65_reset),
    .io_in_a(FP_adder_13ccs_65_io_in_a),
    .io_in_b(FP_adder_13ccs_65_io_in_b),
    .io_out_s(FP_adder_13ccs_65_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_66 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_66_clock),
    .reset(FP_adder_13ccs_66_reset),
    .io_in_a(FP_adder_13ccs_66_io_in_a),
    .io_in_b(FP_adder_13ccs_66_io_in_b),
    .io_out_s(FP_adder_13ccs_66_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_67 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_67_clock),
    .reset(FP_adder_13ccs_67_reset),
    .io_in_a(FP_adder_13ccs_67_io_in_a),
    .io_in_b(FP_adder_13ccs_67_io_in_b),
    .io_out_s(FP_adder_13ccs_67_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_68 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_68_clock),
    .reset(FP_adder_13ccs_68_reset),
    .io_in_a(FP_adder_13ccs_68_io_in_a),
    .io_in_b(FP_adder_13ccs_68_io_in_b),
    .io_out_s(FP_adder_13ccs_68_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_69 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_69_clock),
    .reset(FP_adder_13ccs_69_reset),
    .io_in_a(FP_adder_13ccs_69_io_in_a),
    .io_in_b(FP_adder_13ccs_69_io_in_b),
    .io_out_s(FP_adder_13ccs_69_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_70 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_70_clock),
    .reset(FP_adder_13ccs_70_reset),
    .io_in_a(FP_adder_13ccs_70_io_in_a),
    .io_in_b(FP_adder_13ccs_70_io_in_b),
    .io_out_s(FP_adder_13ccs_70_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_71 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_71_clock),
    .reset(FP_adder_13ccs_71_reset),
    .io_in_a(FP_adder_13ccs_71_io_in_a),
    .io_in_b(FP_adder_13ccs_71_io_in_b),
    .io_out_s(FP_adder_13ccs_71_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_72 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_72_clock),
    .reset(FP_adder_13ccs_72_reset),
    .io_in_a(FP_adder_13ccs_72_io_in_a),
    .io_in_b(FP_adder_13ccs_72_io_in_b),
    .io_out_s(FP_adder_13ccs_72_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_73 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_73_clock),
    .reset(FP_adder_13ccs_73_reset),
    .io_in_a(FP_adder_13ccs_73_io_in_a),
    .io_in_b(FP_adder_13ccs_73_io_in_b),
    .io_out_s(FP_adder_13ccs_73_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_74 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_74_clock),
    .reset(FP_adder_13ccs_74_reset),
    .io_in_a(FP_adder_13ccs_74_io_in_a),
    .io_in_b(FP_adder_13ccs_74_io_in_b),
    .io_out_s(FP_adder_13ccs_74_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_75 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_75_clock),
    .reset(FP_adder_13ccs_75_reset),
    .io_in_a(FP_adder_13ccs_75_io_in_a),
    .io_in_b(FP_adder_13ccs_75_io_in_b),
    .io_out_s(FP_adder_13ccs_75_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_76 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_76_clock),
    .reset(FP_adder_13ccs_76_reset),
    .io_in_a(FP_adder_13ccs_76_io_in_a),
    .io_in_b(FP_adder_13ccs_76_io_in_b),
    .io_out_s(FP_adder_13ccs_76_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_77 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_77_clock),
    .reset(FP_adder_13ccs_77_reset),
    .io_in_a(FP_adder_13ccs_77_io_in_a),
    .io_in_b(FP_adder_13ccs_77_io_in_b),
    .io_out_s(FP_adder_13ccs_77_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_78 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_78_clock),
    .reset(FP_adder_13ccs_78_reset),
    .io_in_a(FP_adder_13ccs_78_io_in_a),
    .io_in_b(FP_adder_13ccs_78_io_in_b),
    .io_out_s(FP_adder_13ccs_78_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_79 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_79_clock),
    .reset(FP_adder_13ccs_79_reset),
    .io_in_a(FP_adder_13ccs_79_io_in_a),
    .io_in_b(FP_adder_13ccs_79_io_in_b),
    .io_out_s(FP_adder_13ccs_79_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_80 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_80_clock),
    .reset(FP_adder_13ccs_80_reset),
    .io_in_a(FP_adder_13ccs_80_io_in_a),
    .io_in_b(FP_adder_13ccs_80_io_in_b),
    .io_out_s(FP_adder_13ccs_80_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_81 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_81_clock),
    .reset(FP_adder_13ccs_81_reset),
    .io_in_a(FP_adder_13ccs_81_io_in_a),
    .io_in_b(FP_adder_13ccs_81_io_in_b),
    .io_out_s(FP_adder_13ccs_81_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_82 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_82_clock),
    .reset(FP_adder_13ccs_82_reset),
    .io_in_a(FP_adder_13ccs_82_io_in_a),
    .io_in_b(FP_adder_13ccs_82_io_in_b),
    .io_out_s(FP_adder_13ccs_82_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_83 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_83_clock),
    .reset(FP_adder_13ccs_83_reset),
    .io_in_a(FP_adder_13ccs_83_io_in_a),
    .io_in_b(FP_adder_13ccs_83_io_in_b),
    .io_out_s(FP_adder_13ccs_83_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_84 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_84_clock),
    .reset(FP_adder_13ccs_84_reset),
    .io_in_a(FP_adder_13ccs_84_io_in_a),
    .io_in_b(FP_adder_13ccs_84_io_in_b),
    .io_out_s(FP_adder_13ccs_84_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_85 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_85_clock),
    .reset(FP_adder_13ccs_85_reset),
    .io_in_a(FP_adder_13ccs_85_io_in_a),
    .io_in_b(FP_adder_13ccs_85_io_in_b),
    .io_out_s(FP_adder_13ccs_85_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_86 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_86_clock),
    .reset(FP_adder_13ccs_86_reset),
    .io_in_a(FP_adder_13ccs_86_io_in_a),
    .io_in_b(FP_adder_13ccs_86_io_in_b),
    .io_out_s(FP_adder_13ccs_86_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_87 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_87_clock),
    .reset(FP_adder_13ccs_87_reset),
    .io_in_a(FP_adder_13ccs_87_io_in_a),
    .io_in_b(FP_adder_13ccs_87_io_in_b),
    .io_out_s(FP_adder_13ccs_87_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_88 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_88_clock),
    .reset(FP_adder_13ccs_88_reset),
    .io_in_a(FP_adder_13ccs_88_io_in_a),
    .io_in_b(FP_adder_13ccs_88_io_in_b),
    .io_out_s(FP_adder_13ccs_88_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_89 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_89_clock),
    .reset(FP_adder_13ccs_89_reset),
    .io_in_a(FP_adder_13ccs_89_io_in_a),
    .io_in_b(FP_adder_13ccs_89_io_in_b),
    .io_out_s(FP_adder_13ccs_89_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_90 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_90_clock),
    .reset(FP_adder_13ccs_90_reset),
    .io_in_a(FP_adder_13ccs_90_io_in_a),
    .io_in_b(FP_adder_13ccs_90_io_in_b),
    .io_out_s(FP_adder_13ccs_90_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_91 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_91_clock),
    .reset(FP_adder_13ccs_91_reset),
    .io_in_a(FP_adder_13ccs_91_io_in_a),
    .io_in_b(FP_adder_13ccs_91_io_in_b),
    .io_out_s(FP_adder_13ccs_91_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_92 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_92_clock),
    .reset(FP_adder_13ccs_92_reset),
    .io_in_a(FP_adder_13ccs_92_io_in_a),
    .io_in_b(FP_adder_13ccs_92_io_in_b),
    .io_out_s(FP_adder_13ccs_92_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_93 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_93_clock),
    .reset(FP_adder_13ccs_93_reset),
    .io_in_a(FP_adder_13ccs_93_io_in_a),
    .io_in_b(FP_adder_13ccs_93_io_in_b),
    .io_out_s(FP_adder_13ccs_93_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_94 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_94_clock),
    .reset(FP_adder_13ccs_94_reset),
    .io_in_a(FP_adder_13ccs_94_io_in_a),
    .io_in_b(FP_adder_13ccs_94_io_in_b),
    .io_out_s(FP_adder_13ccs_94_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_95 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_95_clock),
    .reset(FP_adder_13ccs_95_reset),
    .io_in_a(FP_adder_13ccs_95_io_in_a),
    .io_in_b(FP_adder_13ccs_95_io_in_b),
    .io_out_s(FP_adder_13ccs_95_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_96 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_96_clock),
    .reset(FP_adder_13ccs_96_reset),
    .io_in_a(FP_adder_13ccs_96_io_in_a),
    .io_in_b(FP_adder_13ccs_96_io_in_b),
    .io_out_s(FP_adder_13ccs_96_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_97 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_97_clock),
    .reset(FP_adder_13ccs_97_reset),
    .io_in_a(FP_adder_13ccs_97_io_in_a),
    .io_in_b(FP_adder_13ccs_97_io_in_b),
    .io_out_s(FP_adder_13ccs_97_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_98 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_98_clock),
    .reset(FP_adder_13ccs_98_reset),
    .io_in_a(FP_adder_13ccs_98_io_in_a),
    .io_in_b(FP_adder_13ccs_98_io_in_b),
    .io_out_s(FP_adder_13ccs_98_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_99 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_99_clock),
    .reset(FP_adder_13ccs_99_reset),
    .io_in_a(FP_adder_13ccs_99_io_in_a),
    .io_in_b(FP_adder_13ccs_99_io_in_b),
    .io_out_s(FP_adder_13ccs_99_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_100 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_100_clock),
    .reset(FP_adder_13ccs_100_reset),
    .io_in_a(FP_adder_13ccs_100_io_in_a),
    .io_in_b(FP_adder_13ccs_100_io_in_b),
    .io_out_s(FP_adder_13ccs_100_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_101 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_101_clock),
    .reset(FP_adder_13ccs_101_reset),
    .io_in_a(FP_adder_13ccs_101_io_in_a),
    .io_in_b(FP_adder_13ccs_101_io_in_b),
    .io_out_s(FP_adder_13ccs_101_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_102 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_102_clock),
    .reset(FP_adder_13ccs_102_reset),
    .io_in_a(FP_adder_13ccs_102_io_in_a),
    .io_in_b(FP_adder_13ccs_102_io_in_b),
    .io_out_s(FP_adder_13ccs_102_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_103 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_103_clock),
    .reset(FP_adder_13ccs_103_reset),
    .io_in_a(FP_adder_13ccs_103_io_in_a),
    .io_in_b(FP_adder_13ccs_103_io_in_b),
    .io_out_s(FP_adder_13ccs_103_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_104 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_104_clock),
    .reset(FP_adder_13ccs_104_reset),
    .io_in_a(FP_adder_13ccs_104_io_in_a),
    .io_in_b(FP_adder_13ccs_104_io_in_b),
    .io_out_s(FP_adder_13ccs_104_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_105 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_105_clock),
    .reset(FP_adder_13ccs_105_reset),
    .io_in_a(FP_adder_13ccs_105_io_in_a),
    .io_in_b(FP_adder_13ccs_105_io_in_b),
    .io_out_s(FP_adder_13ccs_105_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_106 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_106_clock),
    .reset(FP_adder_13ccs_106_reset),
    .io_in_a(FP_adder_13ccs_106_io_in_a),
    .io_in_b(FP_adder_13ccs_106_io_in_b),
    .io_out_s(FP_adder_13ccs_106_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_107 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_107_clock),
    .reset(FP_adder_13ccs_107_reset),
    .io_in_a(FP_adder_13ccs_107_io_in_a),
    .io_in_b(FP_adder_13ccs_107_io_in_b),
    .io_out_s(FP_adder_13ccs_107_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_108 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_108_clock),
    .reset(FP_adder_13ccs_108_reset),
    .io_in_a(FP_adder_13ccs_108_io_in_a),
    .io_in_b(FP_adder_13ccs_108_io_in_b),
    .io_out_s(FP_adder_13ccs_108_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_109 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_109_clock),
    .reset(FP_adder_13ccs_109_reset),
    .io_in_a(FP_adder_13ccs_109_io_in_a),
    .io_in_b(FP_adder_13ccs_109_io_in_b),
    .io_out_s(FP_adder_13ccs_109_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_110 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_110_clock),
    .reset(FP_adder_13ccs_110_reset),
    .io_in_a(FP_adder_13ccs_110_io_in_a),
    .io_in_b(FP_adder_13ccs_110_io_in_b),
    .io_out_s(FP_adder_13ccs_110_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_111 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_111_clock),
    .reset(FP_adder_13ccs_111_reset),
    .io_in_a(FP_adder_13ccs_111_io_in_a),
    .io_in_b(FP_adder_13ccs_111_io_in_b),
    .io_out_s(FP_adder_13ccs_111_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_112 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_112_clock),
    .reset(FP_adder_13ccs_112_reset),
    .io_in_a(FP_adder_13ccs_112_io_in_a),
    .io_in_b(FP_adder_13ccs_112_io_in_b),
    .io_out_s(FP_adder_13ccs_112_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_113 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_113_clock),
    .reset(FP_adder_13ccs_113_reset),
    .io_in_a(FP_adder_13ccs_113_io_in_a),
    .io_in_b(FP_adder_13ccs_113_io_in_b),
    .io_out_s(FP_adder_13ccs_113_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_114 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_114_clock),
    .reset(FP_adder_13ccs_114_reset),
    .io_in_a(FP_adder_13ccs_114_io_in_a),
    .io_in_b(FP_adder_13ccs_114_io_in_b),
    .io_out_s(FP_adder_13ccs_114_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_115 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_115_clock),
    .reset(FP_adder_13ccs_115_reset),
    .io_in_a(FP_adder_13ccs_115_io_in_a),
    .io_in_b(FP_adder_13ccs_115_io_in_b),
    .io_out_s(FP_adder_13ccs_115_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_116 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_116_clock),
    .reset(FP_adder_13ccs_116_reset),
    .io_in_a(FP_adder_13ccs_116_io_in_a),
    .io_in_b(FP_adder_13ccs_116_io_in_b),
    .io_out_s(FP_adder_13ccs_116_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_117 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_117_clock),
    .reset(FP_adder_13ccs_117_reset),
    .io_in_a(FP_adder_13ccs_117_io_in_a),
    .io_in_b(FP_adder_13ccs_117_io_in_b),
    .io_out_s(FP_adder_13ccs_117_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_118 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_118_clock),
    .reset(FP_adder_13ccs_118_reset),
    .io_in_a(FP_adder_13ccs_118_io_in_a),
    .io_in_b(FP_adder_13ccs_118_io_in_b),
    .io_out_s(FP_adder_13ccs_118_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_119 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_119_clock),
    .reset(FP_adder_13ccs_119_reset),
    .io_in_a(FP_adder_13ccs_119_io_in_a),
    .io_in_b(FP_adder_13ccs_119_io_in_b),
    .io_out_s(FP_adder_13ccs_119_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_120 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_120_clock),
    .reset(FP_adder_13ccs_120_reset),
    .io_in_a(FP_adder_13ccs_120_io_in_a),
    .io_in_b(FP_adder_13ccs_120_io_in_b),
    .io_out_s(FP_adder_13ccs_120_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_121 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_121_clock),
    .reset(FP_adder_13ccs_121_reset),
    .io_in_a(FP_adder_13ccs_121_io_in_a),
    .io_in_b(FP_adder_13ccs_121_io_in_b),
    .io_out_s(FP_adder_13ccs_121_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_122 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_122_clock),
    .reset(FP_adder_13ccs_122_reset),
    .io_in_a(FP_adder_13ccs_122_io_in_a),
    .io_in_b(FP_adder_13ccs_122_io_in_b),
    .io_out_s(FP_adder_13ccs_122_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_123 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_123_clock),
    .reset(FP_adder_13ccs_123_reset),
    .io_in_a(FP_adder_13ccs_123_io_in_a),
    .io_in_b(FP_adder_13ccs_123_io_in_b),
    .io_out_s(FP_adder_13ccs_123_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_124 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_124_clock),
    .reset(FP_adder_13ccs_124_reset),
    .io_in_a(FP_adder_13ccs_124_io_in_a),
    .io_in_b(FP_adder_13ccs_124_io_in_b),
    .io_out_s(FP_adder_13ccs_124_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_125 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_125_clock),
    .reset(FP_adder_13ccs_125_reset),
    .io_in_a(FP_adder_13ccs_125_io_in_a),
    .io_in_b(FP_adder_13ccs_125_io_in_b),
    .io_out_s(FP_adder_13ccs_125_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_126 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_126_clock),
    .reset(FP_adder_13ccs_126_reset),
    .io_in_a(FP_adder_13ccs_126_io_in_a),
    .io_in_b(FP_adder_13ccs_126_io_in_b),
    .io_out_s(FP_adder_13ccs_126_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_127 ( // @[FloatingPointDesigns.scala 2488:25]
    .clock(FP_adder_13ccs_127_clock),
    .reset(FP_adder_13ccs_127_reset),
    .io_in_a(FP_adder_13ccs_127_io_in_a),
    .io_in_b(FP_adder_13ccs_127_io_in_b),
    .io_out_s(FP_adder_13ccs_127_io_out_s)
  );
  FPReg FPReg ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_clock),
    .reset(FPReg_reset),
    .io_in(FPReg_io_in),
    .io_out(FPReg_io_out)
  );
  FPReg FPReg_1 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_1_clock),
    .reset(FPReg_1_reset),
    .io_in(FPReg_1_io_in),
    .io_out(FPReg_1_io_out)
  );
  FPReg FPReg_2 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_2_clock),
    .reset(FPReg_2_reset),
    .io_in(FPReg_2_io_in),
    .io_out(FPReg_2_io_out)
  );
  FPReg FPReg_3 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_3_clock),
    .reset(FPReg_3_reset),
    .io_in(FPReg_3_io_in),
    .io_out(FPReg_3_io_out)
  );
  FPReg FPReg_4 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_4_clock),
    .reset(FPReg_4_reset),
    .io_in(FPReg_4_io_in),
    .io_out(FPReg_4_io_out)
  );
  FPReg FPReg_5 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_5_clock),
    .reset(FPReg_5_reset),
    .io_in(FPReg_5_io_in),
    .io_out(FPReg_5_io_out)
  );
  FPReg FPReg_6 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_6_clock),
    .reset(FPReg_6_reset),
    .io_in(FPReg_6_io_in),
    .io_out(FPReg_6_io_out)
  );
  FPReg FPReg_7 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_7_clock),
    .reset(FPReg_7_reset),
    .io_in(FPReg_7_io_in),
    .io_out(FPReg_7_io_out)
  );
  FPReg FPReg_8 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_8_clock),
    .reset(FPReg_8_reset),
    .io_in(FPReg_8_io_in),
    .io_out(FPReg_8_io_out)
  );
  FPReg FPReg_9 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_9_clock),
    .reset(FPReg_9_reset),
    .io_in(FPReg_9_io_in),
    .io_out(FPReg_9_io_out)
  );
  FPReg FPReg_10 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_10_clock),
    .reset(FPReg_10_reset),
    .io_in(FPReg_10_io_in),
    .io_out(FPReg_10_io_out)
  );
  FPReg FPReg_11 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_11_clock),
    .reset(FPReg_11_reset),
    .io_in(FPReg_11_io_in),
    .io_out(FPReg_11_io_out)
  );
  FPReg FPReg_12 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_12_clock),
    .reset(FPReg_12_reset),
    .io_in(FPReg_12_io_in),
    .io_out(FPReg_12_io_out)
  );
  FPReg FPReg_13 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_13_clock),
    .reset(FPReg_13_reset),
    .io_in(FPReg_13_io_in),
    .io_out(FPReg_13_io_out)
  );
  FPReg FPReg_14 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_14_clock),
    .reset(FPReg_14_reset),
    .io_in(FPReg_14_io_in),
    .io_out(FPReg_14_io_out)
  );
  FPReg FPReg_15 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_15_clock),
    .reset(FPReg_15_reset),
    .io_in(FPReg_15_io_in),
    .io_out(FPReg_15_io_out)
  );
  FPReg FPReg_16 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_16_clock),
    .reset(FPReg_16_reset),
    .io_in(FPReg_16_io_in),
    .io_out(FPReg_16_io_out)
  );
  FPReg FPReg_17 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_17_clock),
    .reset(FPReg_17_reset),
    .io_in(FPReg_17_io_in),
    .io_out(FPReg_17_io_out)
  );
  FPReg FPReg_18 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_18_clock),
    .reset(FPReg_18_reset),
    .io_in(FPReg_18_io_in),
    .io_out(FPReg_18_io_out)
  );
  FPReg FPReg_19 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_19_clock),
    .reset(FPReg_19_reset),
    .io_in(FPReg_19_io_in),
    .io_out(FPReg_19_io_out)
  );
  FPReg FPReg_20 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_20_clock),
    .reset(FPReg_20_reset),
    .io_in(FPReg_20_io_in),
    .io_out(FPReg_20_io_out)
  );
  FPReg FPReg_21 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_21_clock),
    .reset(FPReg_21_reset),
    .io_in(FPReg_21_io_in),
    .io_out(FPReg_21_io_out)
  );
  FPReg FPReg_22 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_22_clock),
    .reset(FPReg_22_reset),
    .io_in(FPReg_22_io_in),
    .io_out(FPReg_22_io_out)
  );
  FPReg FPReg_23 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_23_clock),
    .reset(FPReg_23_reset),
    .io_in(FPReg_23_io_in),
    .io_out(FPReg_23_io_out)
  );
  FPReg FPReg_24 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_24_clock),
    .reset(FPReg_24_reset),
    .io_in(FPReg_24_io_in),
    .io_out(FPReg_24_io_out)
  );
  FPReg FPReg_25 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_25_clock),
    .reset(FPReg_25_reset),
    .io_in(FPReg_25_io_in),
    .io_out(FPReg_25_io_out)
  );
  FPReg FPReg_26 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_26_clock),
    .reset(FPReg_26_reset),
    .io_in(FPReg_26_io_in),
    .io_out(FPReg_26_io_out)
  );
  FPReg FPReg_27 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_27_clock),
    .reset(FPReg_27_reset),
    .io_in(FPReg_27_io_in),
    .io_out(FPReg_27_io_out)
  );
  FPReg FPReg_28 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_28_clock),
    .reset(FPReg_28_reset),
    .io_in(FPReg_28_io_in),
    .io_out(FPReg_28_io_out)
  );
  FPReg FPReg_29 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_29_clock),
    .reset(FPReg_29_reset),
    .io_in(FPReg_29_io_in),
    .io_out(FPReg_29_io_out)
  );
  FPReg FPReg_30 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_30_clock),
    .reset(FPReg_30_reset),
    .io_in(FPReg_30_io_in),
    .io_out(FPReg_30_io_out)
  );
  FPReg FPReg_31 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_31_clock),
    .reset(FPReg_31_reset),
    .io_in(FPReg_31_io_in),
    .io_out(FPReg_31_io_out)
  );
  FPReg FPReg_32 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_32_clock),
    .reset(FPReg_32_reset),
    .io_in(FPReg_32_io_in),
    .io_out(FPReg_32_io_out)
  );
  FPReg FPReg_33 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_33_clock),
    .reset(FPReg_33_reset),
    .io_in(FPReg_33_io_in),
    .io_out(FPReg_33_io_out)
  );
  FPReg FPReg_34 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_34_clock),
    .reset(FPReg_34_reset),
    .io_in(FPReg_34_io_in),
    .io_out(FPReg_34_io_out)
  );
  FPReg FPReg_35 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_35_clock),
    .reset(FPReg_35_reset),
    .io_in(FPReg_35_io_in),
    .io_out(FPReg_35_io_out)
  );
  FPReg FPReg_36 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_36_clock),
    .reset(FPReg_36_reset),
    .io_in(FPReg_36_io_in),
    .io_out(FPReg_36_io_out)
  );
  FPReg FPReg_37 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_37_clock),
    .reset(FPReg_37_reset),
    .io_in(FPReg_37_io_in),
    .io_out(FPReg_37_io_out)
  );
  FPReg FPReg_38 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_38_clock),
    .reset(FPReg_38_reset),
    .io_in(FPReg_38_io_in),
    .io_out(FPReg_38_io_out)
  );
  FPReg FPReg_39 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_39_clock),
    .reset(FPReg_39_reset),
    .io_in(FPReg_39_io_in),
    .io_out(FPReg_39_io_out)
  );
  FPReg FPReg_40 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_40_clock),
    .reset(FPReg_40_reset),
    .io_in(FPReg_40_io_in),
    .io_out(FPReg_40_io_out)
  );
  FPReg FPReg_41 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_41_clock),
    .reset(FPReg_41_reset),
    .io_in(FPReg_41_io_in),
    .io_out(FPReg_41_io_out)
  );
  FPReg FPReg_42 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_42_clock),
    .reset(FPReg_42_reset),
    .io_in(FPReg_42_io_in),
    .io_out(FPReg_42_io_out)
  );
  FPReg FPReg_43 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_43_clock),
    .reset(FPReg_43_reset),
    .io_in(FPReg_43_io_in),
    .io_out(FPReg_43_io_out)
  );
  FPReg FPReg_44 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_44_clock),
    .reset(FPReg_44_reset),
    .io_in(FPReg_44_io_in),
    .io_out(FPReg_44_io_out)
  );
  FPReg FPReg_45 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_45_clock),
    .reset(FPReg_45_reset),
    .io_in(FPReg_45_io_in),
    .io_out(FPReg_45_io_out)
  );
  FPReg FPReg_46 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_46_clock),
    .reset(FPReg_46_reset),
    .io_in(FPReg_46_io_in),
    .io_out(FPReg_46_io_out)
  );
  FPReg FPReg_47 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_47_clock),
    .reset(FPReg_47_reset),
    .io_in(FPReg_47_io_in),
    .io_out(FPReg_47_io_out)
  );
  FPReg FPReg_48 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_48_clock),
    .reset(FPReg_48_reset),
    .io_in(FPReg_48_io_in),
    .io_out(FPReg_48_io_out)
  );
  FPReg FPReg_49 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_49_clock),
    .reset(FPReg_49_reset),
    .io_in(FPReg_49_io_in),
    .io_out(FPReg_49_io_out)
  );
  FPReg FPReg_50 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_50_clock),
    .reset(FPReg_50_reset),
    .io_in(FPReg_50_io_in),
    .io_out(FPReg_50_io_out)
  );
  FPReg FPReg_51 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_51_clock),
    .reset(FPReg_51_reset),
    .io_in(FPReg_51_io_in),
    .io_out(FPReg_51_io_out)
  );
  FPReg FPReg_52 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_52_clock),
    .reset(FPReg_52_reset),
    .io_in(FPReg_52_io_in),
    .io_out(FPReg_52_io_out)
  );
  FPReg FPReg_53 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_53_clock),
    .reset(FPReg_53_reset),
    .io_in(FPReg_53_io_in),
    .io_out(FPReg_53_io_out)
  );
  FPReg FPReg_54 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_54_clock),
    .reset(FPReg_54_reset),
    .io_in(FPReg_54_io_in),
    .io_out(FPReg_54_io_out)
  );
  FPReg FPReg_55 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_55_clock),
    .reset(FPReg_55_reset),
    .io_in(FPReg_55_io_in),
    .io_out(FPReg_55_io_out)
  );
  FPReg FPReg_56 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_56_clock),
    .reset(FPReg_56_reset),
    .io_in(FPReg_56_io_in),
    .io_out(FPReg_56_io_out)
  );
  FPReg FPReg_57 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_57_clock),
    .reset(FPReg_57_reset),
    .io_in(FPReg_57_io_in),
    .io_out(FPReg_57_io_out)
  );
  FPReg FPReg_58 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_58_clock),
    .reset(FPReg_58_reset),
    .io_in(FPReg_58_io_in),
    .io_out(FPReg_58_io_out)
  );
  FPReg FPReg_59 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_59_clock),
    .reset(FPReg_59_reset),
    .io_in(FPReg_59_io_in),
    .io_out(FPReg_59_io_out)
  );
  FPReg FPReg_60 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_60_clock),
    .reset(FPReg_60_reset),
    .io_in(FPReg_60_io_in),
    .io_out(FPReg_60_io_out)
  );
  FPReg FPReg_61 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_61_clock),
    .reset(FPReg_61_reset),
    .io_in(FPReg_61_io_in),
    .io_out(FPReg_61_io_out)
  );
  FPReg FPReg_62 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_62_clock),
    .reset(FPReg_62_reset),
    .io_in(FPReg_62_io_in),
    .io_out(FPReg_62_io_out)
  );
  FPReg FPReg_63 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_63_clock),
    .reset(FPReg_63_reset),
    .io_in(FPReg_63_io_in),
    .io_out(FPReg_63_io_out)
  );
  FPReg FPReg_64 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_64_clock),
    .reset(FPReg_64_reset),
    .io_in(FPReg_64_io_in),
    .io_out(FPReg_64_io_out)
  );
  FPReg FPReg_65 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_65_clock),
    .reset(FPReg_65_reset),
    .io_in(FPReg_65_io_in),
    .io_out(FPReg_65_io_out)
  );
  FPReg FPReg_66 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_66_clock),
    .reset(FPReg_66_reset),
    .io_in(FPReg_66_io_in),
    .io_out(FPReg_66_io_out)
  );
  FPReg FPReg_67 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_67_clock),
    .reset(FPReg_67_reset),
    .io_in(FPReg_67_io_in),
    .io_out(FPReg_67_io_out)
  );
  FPReg FPReg_68 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_68_clock),
    .reset(FPReg_68_reset),
    .io_in(FPReg_68_io_in),
    .io_out(FPReg_68_io_out)
  );
  FPReg FPReg_69 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_69_clock),
    .reset(FPReg_69_reset),
    .io_in(FPReg_69_io_in),
    .io_out(FPReg_69_io_out)
  );
  FPReg FPReg_70 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_70_clock),
    .reset(FPReg_70_reset),
    .io_in(FPReg_70_io_in),
    .io_out(FPReg_70_io_out)
  );
  FPReg FPReg_71 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_71_clock),
    .reset(FPReg_71_reset),
    .io_in(FPReg_71_io_in),
    .io_out(FPReg_71_io_out)
  );
  FPReg FPReg_72 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_72_clock),
    .reset(FPReg_72_reset),
    .io_in(FPReg_72_io_in),
    .io_out(FPReg_72_io_out)
  );
  FPReg FPReg_73 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_73_clock),
    .reset(FPReg_73_reset),
    .io_in(FPReg_73_io_in),
    .io_out(FPReg_73_io_out)
  );
  FPReg FPReg_74 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_74_clock),
    .reset(FPReg_74_reset),
    .io_in(FPReg_74_io_in),
    .io_out(FPReg_74_io_out)
  );
  FPReg FPReg_75 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_75_clock),
    .reset(FPReg_75_reset),
    .io_in(FPReg_75_io_in),
    .io_out(FPReg_75_io_out)
  );
  FPReg FPReg_76 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_76_clock),
    .reset(FPReg_76_reset),
    .io_in(FPReg_76_io_in),
    .io_out(FPReg_76_io_out)
  );
  FPReg FPReg_77 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_77_clock),
    .reset(FPReg_77_reset),
    .io_in(FPReg_77_io_in),
    .io_out(FPReg_77_io_out)
  );
  FPReg FPReg_78 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_78_clock),
    .reset(FPReg_78_reset),
    .io_in(FPReg_78_io_in),
    .io_out(FPReg_78_io_out)
  );
  FPReg FPReg_79 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_79_clock),
    .reset(FPReg_79_reset),
    .io_in(FPReg_79_io_in),
    .io_out(FPReg_79_io_out)
  );
  FPReg FPReg_80 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_80_clock),
    .reset(FPReg_80_reset),
    .io_in(FPReg_80_io_in),
    .io_out(FPReg_80_io_out)
  );
  FPReg FPReg_81 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_81_clock),
    .reset(FPReg_81_reset),
    .io_in(FPReg_81_io_in),
    .io_out(FPReg_81_io_out)
  );
  FPReg FPReg_82 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_82_clock),
    .reset(FPReg_82_reset),
    .io_in(FPReg_82_io_in),
    .io_out(FPReg_82_io_out)
  );
  FPReg FPReg_83 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_83_clock),
    .reset(FPReg_83_reset),
    .io_in(FPReg_83_io_in),
    .io_out(FPReg_83_io_out)
  );
  FPReg FPReg_84 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_84_clock),
    .reset(FPReg_84_reset),
    .io_in(FPReg_84_io_in),
    .io_out(FPReg_84_io_out)
  );
  FPReg FPReg_85 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_85_clock),
    .reset(FPReg_85_reset),
    .io_in(FPReg_85_io_in),
    .io_out(FPReg_85_io_out)
  );
  FPReg FPReg_86 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_86_clock),
    .reset(FPReg_86_reset),
    .io_in(FPReg_86_io_in),
    .io_out(FPReg_86_io_out)
  );
  FPReg FPReg_87 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_87_clock),
    .reset(FPReg_87_reset),
    .io_in(FPReg_87_io_in),
    .io_out(FPReg_87_io_out)
  );
  FPReg FPReg_88 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_88_clock),
    .reset(FPReg_88_reset),
    .io_in(FPReg_88_io_in),
    .io_out(FPReg_88_io_out)
  );
  FPReg FPReg_89 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_89_clock),
    .reset(FPReg_89_reset),
    .io_in(FPReg_89_io_in),
    .io_out(FPReg_89_io_out)
  );
  FPReg FPReg_90 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_90_clock),
    .reset(FPReg_90_reset),
    .io_in(FPReg_90_io_in),
    .io_out(FPReg_90_io_out)
  );
  FPReg FPReg_91 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_91_clock),
    .reset(FPReg_91_reset),
    .io_in(FPReg_91_io_in),
    .io_out(FPReg_91_io_out)
  );
  FPReg FPReg_92 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_92_clock),
    .reset(FPReg_92_reset),
    .io_in(FPReg_92_io_in),
    .io_out(FPReg_92_io_out)
  );
  FPReg FPReg_93 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_93_clock),
    .reset(FPReg_93_reset),
    .io_in(FPReg_93_io_in),
    .io_out(FPReg_93_io_out)
  );
  FPReg FPReg_94 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_94_clock),
    .reset(FPReg_94_reset),
    .io_in(FPReg_94_io_in),
    .io_out(FPReg_94_io_out)
  );
  FPReg FPReg_95 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_95_clock),
    .reset(FPReg_95_reset),
    .io_in(FPReg_95_io_in),
    .io_out(FPReg_95_io_out)
  );
  FPReg FPReg_96 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_96_clock),
    .reset(FPReg_96_reset),
    .io_in(FPReg_96_io_in),
    .io_out(FPReg_96_io_out)
  );
  FPReg FPReg_97 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_97_clock),
    .reset(FPReg_97_reset),
    .io_in(FPReg_97_io_in),
    .io_out(FPReg_97_io_out)
  );
  FPReg FPReg_98 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_98_clock),
    .reset(FPReg_98_reset),
    .io_in(FPReg_98_io_in),
    .io_out(FPReg_98_io_out)
  );
  FPReg FPReg_99 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_99_clock),
    .reset(FPReg_99_reset),
    .io_in(FPReg_99_io_in),
    .io_out(FPReg_99_io_out)
  );
  FPReg FPReg_100 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_100_clock),
    .reset(FPReg_100_reset),
    .io_in(FPReg_100_io_in),
    .io_out(FPReg_100_io_out)
  );
  FPReg FPReg_101 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_101_clock),
    .reset(FPReg_101_reset),
    .io_in(FPReg_101_io_in),
    .io_out(FPReg_101_io_out)
  );
  FPReg FPReg_102 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_102_clock),
    .reset(FPReg_102_reset),
    .io_in(FPReg_102_io_in),
    .io_out(FPReg_102_io_out)
  );
  FPReg FPReg_103 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_103_clock),
    .reset(FPReg_103_reset),
    .io_in(FPReg_103_io_in),
    .io_out(FPReg_103_io_out)
  );
  FPReg FPReg_104 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_104_clock),
    .reset(FPReg_104_reset),
    .io_in(FPReg_104_io_in),
    .io_out(FPReg_104_io_out)
  );
  FPReg FPReg_105 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_105_clock),
    .reset(FPReg_105_reset),
    .io_in(FPReg_105_io_in),
    .io_out(FPReg_105_io_out)
  );
  FPReg FPReg_106 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_106_clock),
    .reset(FPReg_106_reset),
    .io_in(FPReg_106_io_in),
    .io_out(FPReg_106_io_out)
  );
  FPReg FPReg_107 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_107_clock),
    .reset(FPReg_107_reset),
    .io_in(FPReg_107_io_in),
    .io_out(FPReg_107_io_out)
  );
  FPReg FPReg_108 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_108_clock),
    .reset(FPReg_108_reset),
    .io_in(FPReg_108_io_in),
    .io_out(FPReg_108_io_out)
  );
  FPReg FPReg_109 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_109_clock),
    .reset(FPReg_109_reset),
    .io_in(FPReg_109_io_in),
    .io_out(FPReg_109_io_out)
  );
  FPReg FPReg_110 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_110_clock),
    .reset(FPReg_110_reset),
    .io_in(FPReg_110_io_in),
    .io_out(FPReg_110_io_out)
  );
  FPReg FPReg_111 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_111_clock),
    .reset(FPReg_111_reset),
    .io_in(FPReg_111_io_in),
    .io_out(FPReg_111_io_out)
  );
  FPReg FPReg_112 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_112_clock),
    .reset(FPReg_112_reset),
    .io_in(FPReg_112_io_in),
    .io_out(FPReg_112_io_out)
  );
  FPReg FPReg_113 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_113_clock),
    .reset(FPReg_113_reset),
    .io_in(FPReg_113_io_in),
    .io_out(FPReg_113_io_out)
  );
  FPReg FPReg_114 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_114_clock),
    .reset(FPReg_114_reset),
    .io_in(FPReg_114_io_in),
    .io_out(FPReg_114_io_out)
  );
  FPReg FPReg_115 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_115_clock),
    .reset(FPReg_115_reset),
    .io_in(FPReg_115_io_in),
    .io_out(FPReg_115_io_out)
  );
  FPReg FPReg_116 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_116_clock),
    .reset(FPReg_116_reset),
    .io_in(FPReg_116_io_in),
    .io_out(FPReg_116_io_out)
  );
  FPReg FPReg_117 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_117_clock),
    .reset(FPReg_117_reset),
    .io_in(FPReg_117_io_in),
    .io_out(FPReg_117_io_out)
  );
  FPReg FPReg_118 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_118_clock),
    .reset(FPReg_118_reset),
    .io_in(FPReg_118_io_in),
    .io_out(FPReg_118_io_out)
  );
  FPReg FPReg_119 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_119_clock),
    .reset(FPReg_119_reset),
    .io_in(FPReg_119_io_in),
    .io_out(FPReg_119_io_out)
  );
  FPReg FPReg_120 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_120_clock),
    .reset(FPReg_120_reset),
    .io_in(FPReg_120_io_in),
    .io_out(FPReg_120_io_out)
  );
  FPReg FPReg_121 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_121_clock),
    .reset(FPReg_121_reset),
    .io_in(FPReg_121_io_in),
    .io_out(FPReg_121_io_out)
  );
  FPReg FPReg_122 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_122_clock),
    .reset(FPReg_122_reset),
    .io_in(FPReg_122_io_in),
    .io_out(FPReg_122_io_out)
  );
  FPReg FPReg_123 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_123_clock),
    .reset(FPReg_123_reset),
    .io_in(FPReg_123_io_in),
    .io_out(FPReg_123_io_out)
  );
  FPReg FPReg_124 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_124_clock),
    .reset(FPReg_124_reset),
    .io_in(FPReg_124_io_in),
    .io_out(FPReg_124_io_out)
  );
  FPReg FPReg_125 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_125_clock),
    .reset(FPReg_125_reset),
    .io_in(FPReg_125_io_in),
    .io_out(FPReg_125_io_out)
  );
  FPReg FPReg_126 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_126_clock),
    .reset(FPReg_126_reset),
    .io_in(FPReg_126_io_in),
    .io_out(FPReg_126_io_out)
  );
  FPReg FPReg_127 ( // @[FloatingPointDesigns.scala 2492:48]
    .clock(FPReg_127_clock),
    .reset(FPReg_127_reset),
    .io_in(FPReg_127_io_in),
    .io_out(FPReg_127_io_out)
  );
  assign io_out_s_0 = FP_adder_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_1 = FP_adder_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_2 = FP_adder_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_3 = FP_adder_13ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_4 = FP_adder_13ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_5 = FP_adder_13ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_6 = FP_adder_13ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_7 = FP_adder_13ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_8 = FP_adder_13ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_9 = FP_adder_13ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_10 = FP_adder_13ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_11 = FP_adder_13ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_12 = FP_adder_13ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_13 = FP_adder_13ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_14 = FP_adder_13ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_15 = FP_adder_13ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_16 = FP_adder_13ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_17 = FP_adder_13ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_18 = FP_adder_13ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_19 = FP_adder_13ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_20 = FP_adder_13ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_21 = FP_adder_13ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_22 = FP_adder_13ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_23 = FP_adder_13ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_24 = FP_adder_13ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_25 = FP_adder_13ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_26 = FP_adder_13ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_27 = FP_adder_13ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_28 = FP_adder_13ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_29 = FP_adder_13ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_30 = FP_adder_13ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_31 = FP_adder_13ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_32 = FP_adder_13ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_33 = FP_adder_13ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_34 = FP_adder_13ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_35 = FP_adder_13ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_36 = FP_adder_13ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_37 = FP_adder_13ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_38 = FP_adder_13ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_39 = FP_adder_13ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_40 = FP_adder_13ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_41 = FP_adder_13ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_42 = FP_adder_13ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_43 = FP_adder_13ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_44 = FP_adder_13ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_45 = FP_adder_13ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_46 = FP_adder_13ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_47 = FP_adder_13ccs_47_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_48 = FP_adder_13ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_49 = FP_adder_13ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_50 = FP_adder_13ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_51 = FP_adder_13ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_52 = FP_adder_13ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_53 = FP_adder_13ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_54 = FP_adder_13ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_55 = FP_adder_13ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_56 = FP_adder_13ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_57 = FP_adder_13ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_58 = FP_adder_13ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_59 = FP_adder_13ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_60 = FP_adder_13ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_61 = FP_adder_13ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_62 = FP_adder_13ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_63 = FP_adder_13ccs_63_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_64 = FP_adder_13ccs_64_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_65 = FP_adder_13ccs_65_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_66 = FP_adder_13ccs_66_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_67 = FP_adder_13ccs_67_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_68 = FP_adder_13ccs_68_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_69 = FP_adder_13ccs_69_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_70 = FP_adder_13ccs_70_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_71 = FP_adder_13ccs_71_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_72 = FP_adder_13ccs_72_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_73 = FP_adder_13ccs_73_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_74 = FP_adder_13ccs_74_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_75 = FP_adder_13ccs_75_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_76 = FP_adder_13ccs_76_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_77 = FP_adder_13ccs_77_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_78 = FP_adder_13ccs_78_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_79 = FP_adder_13ccs_79_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_80 = FP_adder_13ccs_80_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_81 = FP_adder_13ccs_81_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_82 = FP_adder_13ccs_82_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_83 = FP_adder_13ccs_83_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_84 = FP_adder_13ccs_84_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_85 = FP_adder_13ccs_85_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_86 = FP_adder_13ccs_86_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_87 = FP_adder_13ccs_87_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_88 = FP_adder_13ccs_88_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_89 = FP_adder_13ccs_89_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_90 = FP_adder_13ccs_90_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_91 = FP_adder_13ccs_91_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_92 = FP_adder_13ccs_92_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_93 = FP_adder_13ccs_93_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_94 = FP_adder_13ccs_94_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_95 = FP_adder_13ccs_95_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_96 = FP_adder_13ccs_96_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_97 = FP_adder_13ccs_97_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_98 = FP_adder_13ccs_98_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_99 = FP_adder_13ccs_99_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_100 = FP_adder_13ccs_100_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_101 = FP_adder_13ccs_101_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_102 = FP_adder_13ccs_102_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_103 = FP_adder_13ccs_103_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_104 = FP_adder_13ccs_104_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_105 = FP_adder_13ccs_105_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_106 = FP_adder_13ccs_106_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_107 = FP_adder_13ccs_107_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_108 = FP_adder_13ccs_108_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_109 = FP_adder_13ccs_109_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_110 = FP_adder_13ccs_110_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_111 = FP_adder_13ccs_111_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_112 = FP_adder_13ccs_112_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_113 = FP_adder_13ccs_113_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_114 = FP_adder_13ccs_114_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_115 = FP_adder_13ccs_115_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_116 = FP_adder_13ccs_116_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_117 = FP_adder_13ccs_117_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_118 = FP_adder_13ccs_118_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_119 = FP_adder_13ccs_119_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_120 = FP_adder_13ccs_120_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_121 = FP_adder_13ccs_121_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_122 = FP_adder_13ccs_122_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_123 = FP_adder_13ccs_123_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_124 = FP_adder_13ccs_124_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_125 = FP_adder_13ccs_125_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_126 = FP_adder_13ccs_126_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign io_out_s_127 = FP_adder_13ccs_127_io_out_s; // @[FloatingPointDesigns.scala 2499:19]
  assign FP_multiplier_10ccs_clock = clock;
  assign FP_multiplier_10ccs_reset = reset;
  assign FP_multiplier_10ccs_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_io_in_b = io_in_b_0; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_1_clock = clock;
  assign FP_multiplier_10ccs_1_reset = reset;
  assign FP_multiplier_10ccs_1_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_1_io_in_b = io_in_b_1; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_2_clock = clock;
  assign FP_multiplier_10ccs_2_reset = reset;
  assign FP_multiplier_10ccs_2_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_2_io_in_b = io_in_b_2; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_3_clock = clock;
  assign FP_multiplier_10ccs_3_reset = reset;
  assign FP_multiplier_10ccs_3_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_3_io_in_b = io_in_b_3; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_4_clock = clock;
  assign FP_multiplier_10ccs_4_reset = reset;
  assign FP_multiplier_10ccs_4_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_4_io_in_b = io_in_b_4; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_5_clock = clock;
  assign FP_multiplier_10ccs_5_reset = reset;
  assign FP_multiplier_10ccs_5_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_5_io_in_b = io_in_b_5; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_6_clock = clock;
  assign FP_multiplier_10ccs_6_reset = reset;
  assign FP_multiplier_10ccs_6_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_6_io_in_b = io_in_b_6; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_7_clock = clock;
  assign FP_multiplier_10ccs_7_reset = reset;
  assign FP_multiplier_10ccs_7_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_7_io_in_b = io_in_b_7; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_8_clock = clock;
  assign FP_multiplier_10ccs_8_reset = reset;
  assign FP_multiplier_10ccs_8_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_8_io_in_b = io_in_b_8; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_9_clock = clock;
  assign FP_multiplier_10ccs_9_reset = reset;
  assign FP_multiplier_10ccs_9_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_9_io_in_b = io_in_b_9; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_10_clock = clock;
  assign FP_multiplier_10ccs_10_reset = reset;
  assign FP_multiplier_10ccs_10_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_10_io_in_b = io_in_b_10; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_11_clock = clock;
  assign FP_multiplier_10ccs_11_reset = reset;
  assign FP_multiplier_10ccs_11_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_11_io_in_b = io_in_b_11; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_12_clock = clock;
  assign FP_multiplier_10ccs_12_reset = reset;
  assign FP_multiplier_10ccs_12_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_12_io_in_b = io_in_b_12; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_13_clock = clock;
  assign FP_multiplier_10ccs_13_reset = reset;
  assign FP_multiplier_10ccs_13_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_13_io_in_b = io_in_b_13; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_14_clock = clock;
  assign FP_multiplier_10ccs_14_reset = reset;
  assign FP_multiplier_10ccs_14_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_14_io_in_b = io_in_b_14; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_15_clock = clock;
  assign FP_multiplier_10ccs_15_reset = reset;
  assign FP_multiplier_10ccs_15_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_15_io_in_b = io_in_b_15; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_16_clock = clock;
  assign FP_multiplier_10ccs_16_reset = reset;
  assign FP_multiplier_10ccs_16_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_16_io_in_b = io_in_b_16; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_17_clock = clock;
  assign FP_multiplier_10ccs_17_reset = reset;
  assign FP_multiplier_10ccs_17_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_17_io_in_b = io_in_b_17; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_18_clock = clock;
  assign FP_multiplier_10ccs_18_reset = reset;
  assign FP_multiplier_10ccs_18_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_18_io_in_b = io_in_b_18; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_19_clock = clock;
  assign FP_multiplier_10ccs_19_reset = reset;
  assign FP_multiplier_10ccs_19_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_19_io_in_b = io_in_b_19; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_20_clock = clock;
  assign FP_multiplier_10ccs_20_reset = reset;
  assign FP_multiplier_10ccs_20_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_20_io_in_b = io_in_b_20; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_21_clock = clock;
  assign FP_multiplier_10ccs_21_reset = reset;
  assign FP_multiplier_10ccs_21_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_21_io_in_b = io_in_b_21; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_22_clock = clock;
  assign FP_multiplier_10ccs_22_reset = reset;
  assign FP_multiplier_10ccs_22_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_22_io_in_b = io_in_b_22; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_23_clock = clock;
  assign FP_multiplier_10ccs_23_reset = reset;
  assign FP_multiplier_10ccs_23_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_23_io_in_b = io_in_b_23; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_24_clock = clock;
  assign FP_multiplier_10ccs_24_reset = reset;
  assign FP_multiplier_10ccs_24_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_24_io_in_b = io_in_b_24; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_25_clock = clock;
  assign FP_multiplier_10ccs_25_reset = reset;
  assign FP_multiplier_10ccs_25_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_25_io_in_b = io_in_b_25; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_26_clock = clock;
  assign FP_multiplier_10ccs_26_reset = reset;
  assign FP_multiplier_10ccs_26_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_26_io_in_b = io_in_b_26; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_27_clock = clock;
  assign FP_multiplier_10ccs_27_reset = reset;
  assign FP_multiplier_10ccs_27_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_27_io_in_b = io_in_b_27; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_28_clock = clock;
  assign FP_multiplier_10ccs_28_reset = reset;
  assign FP_multiplier_10ccs_28_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_28_io_in_b = io_in_b_28; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_29_clock = clock;
  assign FP_multiplier_10ccs_29_reset = reset;
  assign FP_multiplier_10ccs_29_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_29_io_in_b = io_in_b_29; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_30_clock = clock;
  assign FP_multiplier_10ccs_30_reset = reset;
  assign FP_multiplier_10ccs_30_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_30_io_in_b = io_in_b_30; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_31_clock = clock;
  assign FP_multiplier_10ccs_31_reset = reset;
  assign FP_multiplier_10ccs_31_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_31_io_in_b = io_in_b_31; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_32_clock = clock;
  assign FP_multiplier_10ccs_32_reset = reset;
  assign FP_multiplier_10ccs_32_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_32_io_in_b = io_in_b_32; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_33_clock = clock;
  assign FP_multiplier_10ccs_33_reset = reset;
  assign FP_multiplier_10ccs_33_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_33_io_in_b = io_in_b_33; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_34_clock = clock;
  assign FP_multiplier_10ccs_34_reset = reset;
  assign FP_multiplier_10ccs_34_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_34_io_in_b = io_in_b_34; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_35_clock = clock;
  assign FP_multiplier_10ccs_35_reset = reset;
  assign FP_multiplier_10ccs_35_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_35_io_in_b = io_in_b_35; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_36_clock = clock;
  assign FP_multiplier_10ccs_36_reset = reset;
  assign FP_multiplier_10ccs_36_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_36_io_in_b = io_in_b_36; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_37_clock = clock;
  assign FP_multiplier_10ccs_37_reset = reset;
  assign FP_multiplier_10ccs_37_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_37_io_in_b = io_in_b_37; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_38_clock = clock;
  assign FP_multiplier_10ccs_38_reset = reset;
  assign FP_multiplier_10ccs_38_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_38_io_in_b = io_in_b_38; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_39_clock = clock;
  assign FP_multiplier_10ccs_39_reset = reset;
  assign FP_multiplier_10ccs_39_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_39_io_in_b = io_in_b_39; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_40_clock = clock;
  assign FP_multiplier_10ccs_40_reset = reset;
  assign FP_multiplier_10ccs_40_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_40_io_in_b = io_in_b_40; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_41_clock = clock;
  assign FP_multiplier_10ccs_41_reset = reset;
  assign FP_multiplier_10ccs_41_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_41_io_in_b = io_in_b_41; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_42_clock = clock;
  assign FP_multiplier_10ccs_42_reset = reset;
  assign FP_multiplier_10ccs_42_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_42_io_in_b = io_in_b_42; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_43_clock = clock;
  assign FP_multiplier_10ccs_43_reset = reset;
  assign FP_multiplier_10ccs_43_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_43_io_in_b = io_in_b_43; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_44_clock = clock;
  assign FP_multiplier_10ccs_44_reset = reset;
  assign FP_multiplier_10ccs_44_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_44_io_in_b = io_in_b_44; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_45_clock = clock;
  assign FP_multiplier_10ccs_45_reset = reset;
  assign FP_multiplier_10ccs_45_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_45_io_in_b = io_in_b_45; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_46_clock = clock;
  assign FP_multiplier_10ccs_46_reset = reset;
  assign FP_multiplier_10ccs_46_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_46_io_in_b = io_in_b_46; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_47_clock = clock;
  assign FP_multiplier_10ccs_47_reset = reset;
  assign FP_multiplier_10ccs_47_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_47_io_in_b = io_in_b_47; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_48_clock = clock;
  assign FP_multiplier_10ccs_48_reset = reset;
  assign FP_multiplier_10ccs_48_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_48_io_in_b = io_in_b_48; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_49_clock = clock;
  assign FP_multiplier_10ccs_49_reset = reset;
  assign FP_multiplier_10ccs_49_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_49_io_in_b = io_in_b_49; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_50_clock = clock;
  assign FP_multiplier_10ccs_50_reset = reset;
  assign FP_multiplier_10ccs_50_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_50_io_in_b = io_in_b_50; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_51_clock = clock;
  assign FP_multiplier_10ccs_51_reset = reset;
  assign FP_multiplier_10ccs_51_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_51_io_in_b = io_in_b_51; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_52_clock = clock;
  assign FP_multiplier_10ccs_52_reset = reset;
  assign FP_multiplier_10ccs_52_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_52_io_in_b = io_in_b_52; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_53_clock = clock;
  assign FP_multiplier_10ccs_53_reset = reset;
  assign FP_multiplier_10ccs_53_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_53_io_in_b = io_in_b_53; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_54_clock = clock;
  assign FP_multiplier_10ccs_54_reset = reset;
  assign FP_multiplier_10ccs_54_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_54_io_in_b = io_in_b_54; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_55_clock = clock;
  assign FP_multiplier_10ccs_55_reset = reset;
  assign FP_multiplier_10ccs_55_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_55_io_in_b = io_in_b_55; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_56_clock = clock;
  assign FP_multiplier_10ccs_56_reset = reset;
  assign FP_multiplier_10ccs_56_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_56_io_in_b = io_in_b_56; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_57_clock = clock;
  assign FP_multiplier_10ccs_57_reset = reset;
  assign FP_multiplier_10ccs_57_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_57_io_in_b = io_in_b_57; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_58_clock = clock;
  assign FP_multiplier_10ccs_58_reset = reset;
  assign FP_multiplier_10ccs_58_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_58_io_in_b = io_in_b_58; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_59_clock = clock;
  assign FP_multiplier_10ccs_59_reset = reset;
  assign FP_multiplier_10ccs_59_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_59_io_in_b = io_in_b_59; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_60_clock = clock;
  assign FP_multiplier_10ccs_60_reset = reset;
  assign FP_multiplier_10ccs_60_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_60_io_in_b = io_in_b_60; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_61_clock = clock;
  assign FP_multiplier_10ccs_61_reset = reset;
  assign FP_multiplier_10ccs_61_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_61_io_in_b = io_in_b_61; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_62_clock = clock;
  assign FP_multiplier_10ccs_62_reset = reset;
  assign FP_multiplier_10ccs_62_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_62_io_in_b = io_in_b_62; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_63_clock = clock;
  assign FP_multiplier_10ccs_63_reset = reset;
  assign FP_multiplier_10ccs_63_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_63_io_in_b = io_in_b_63; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_64_clock = clock;
  assign FP_multiplier_10ccs_64_reset = reset;
  assign FP_multiplier_10ccs_64_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_64_io_in_b = io_in_b_64; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_65_clock = clock;
  assign FP_multiplier_10ccs_65_reset = reset;
  assign FP_multiplier_10ccs_65_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_65_io_in_b = io_in_b_65; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_66_clock = clock;
  assign FP_multiplier_10ccs_66_reset = reset;
  assign FP_multiplier_10ccs_66_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_66_io_in_b = io_in_b_66; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_67_clock = clock;
  assign FP_multiplier_10ccs_67_reset = reset;
  assign FP_multiplier_10ccs_67_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_67_io_in_b = io_in_b_67; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_68_clock = clock;
  assign FP_multiplier_10ccs_68_reset = reset;
  assign FP_multiplier_10ccs_68_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_68_io_in_b = io_in_b_68; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_69_clock = clock;
  assign FP_multiplier_10ccs_69_reset = reset;
  assign FP_multiplier_10ccs_69_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_69_io_in_b = io_in_b_69; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_70_clock = clock;
  assign FP_multiplier_10ccs_70_reset = reset;
  assign FP_multiplier_10ccs_70_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_70_io_in_b = io_in_b_70; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_71_clock = clock;
  assign FP_multiplier_10ccs_71_reset = reset;
  assign FP_multiplier_10ccs_71_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_71_io_in_b = io_in_b_71; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_72_clock = clock;
  assign FP_multiplier_10ccs_72_reset = reset;
  assign FP_multiplier_10ccs_72_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_72_io_in_b = io_in_b_72; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_73_clock = clock;
  assign FP_multiplier_10ccs_73_reset = reset;
  assign FP_multiplier_10ccs_73_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_73_io_in_b = io_in_b_73; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_74_clock = clock;
  assign FP_multiplier_10ccs_74_reset = reset;
  assign FP_multiplier_10ccs_74_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_74_io_in_b = io_in_b_74; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_75_clock = clock;
  assign FP_multiplier_10ccs_75_reset = reset;
  assign FP_multiplier_10ccs_75_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_75_io_in_b = io_in_b_75; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_76_clock = clock;
  assign FP_multiplier_10ccs_76_reset = reset;
  assign FP_multiplier_10ccs_76_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_76_io_in_b = io_in_b_76; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_77_clock = clock;
  assign FP_multiplier_10ccs_77_reset = reset;
  assign FP_multiplier_10ccs_77_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_77_io_in_b = io_in_b_77; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_78_clock = clock;
  assign FP_multiplier_10ccs_78_reset = reset;
  assign FP_multiplier_10ccs_78_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_78_io_in_b = io_in_b_78; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_79_clock = clock;
  assign FP_multiplier_10ccs_79_reset = reset;
  assign FP_multiplier_10ccs_79_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_79_io_in_b = io_in_b_79; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_80_clock = clock;
  assign FP_multiplier_10ccs_80_reset = reset;
  assign FP_multiplier_10ccs_80_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_80_io_in_b = io_in_b_80; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_81_clock = clock;
  assign FP_multiplier_10ccs_81_reset = reset;
  assign FP_multiplier_10ccs_81_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_81_io_in_b = io_in_b_81; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_82_clock = clock;
  assign FP_multiplier_10ccs_82_reset = reset;
  assign FP_multiplier_10ccs_82_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_82_io_in_b = io_in_b_82; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_83_clock = clock;
  assign FP_multiplier_10ccs_83_reset = reset;
  assign FP_multiplier_10ccs_83_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_83_io_in_b = io_in_b_83; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_84_clock = clock;
  assign FP_multiplier_10ccs_84_reset = reset;
  assign FP_multiplier_10ccs_84_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_84_io_in_b = io_in_b_84; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_85_clock = clock;
  assign FP_multiplier_10ccs_85_reset = reset;
  assign FP_multiplier_10ccs_85_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_85_io_in_b = io_in_b_85; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_86_clock = clock;
  assign FP_multiplier_10ccs_86_reset = reset;
  assign FP_multiplier_10ccs_86_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_86_io_in_b = io_in_b_86; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_87_clock = clock;
  assign FP_multiplier_10ccs_87_reset = reset;
  assign FP_multiplier_10ccs_87_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_87_io_in_b = io_in_b_87; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_88_clock = clock;
  assign FP_multiplier_10ccs_88_reset = reset;
  assign FP_multiplier_10ccs_88_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_88_io_in_b = io_in_b_88; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_89_clock = clock;
  assign FP_multiplier_10ccs_89_reset = reset;
  assign FP_multiplier_10ccs_89_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_89_io_in_b = io_in_b_89; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_90_clock = clock;
  assign FP_multiplier_10ccs_90_reset = reset;
  assign FP_multiplier_10ccs_90_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_90_io_in_b = io_in_b_90; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_91_clock = clock;
  assign FP_multiplier_10ccs_91_reset = reset;
  assign FP_multiplier_10ccs_91_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_91_io_in_b = io_in_b_91; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_92_clock = clock;
  assign FP_multiplier_10ccs_92_reset = reset;
  assign FP_multiplier_10ccs_92_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_92_io_in_b = io_in_b_92; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_93_clock = clock;
  assign FP_multiplier_10ccs_93_reset = reset;
  assign FP_multiplier_10ccs_93_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_93_io_in_b = io_in_b_93; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_94_clock = clock;
  assign FP_multiplier_10ccs_94_reset = reset;
  assign FP_multiplier_10ccs_94_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_94_io_in_b = io_in_b_94; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_95_clock = clock;
  assign FP_multiplier_10ccs_95_reset = reset;
  assign FP_multiplier_10ccs_95_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_95_io_in_b = io_in_b_95; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_96_clock = clock;
  assign FP_multiplier_10ccs_96_reset = reset;
  assign FP_multiplier_10ccs_96_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_96_io_in_b = io_in_b_96; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_97_clock = clock;
  assign FP_multiplier_10ccs_97_reset = reset;
  assign FP_multiplier_10ccs_97_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_97_io_in_b = io_in_b_97; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_98_clock = clock;
  assign FP_multiplier_10ccs_98_reset = reset;
  assign FP_multiplier_10ccs_98_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_98_io_in_b = io_in_b_98; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_99_clock = clock;
  assign FP_multiplier_10ccs_99_reset = reset;
  assign FP_multiplier_10ccs_99_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_99_io_in_b = io_in_b_99; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_100_clock = clock;
  assign FP_multiplier_10ccs_100_reset = reset;
  assign FP_multiplier_10ccs_100_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_100_io_in_b = io_in_b_100; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_101_clock = clock;
  assign FP_multiplier_10ccs_101_reset = reset;
  assign FP_multiplier_10ccs_101_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_101_io_in_b = io_in_b_101; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_102_clock = clock;
  assign FP_multiplier_10ccs_102_reset = reset;
  assign FP_multiplier_10ccs_102_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_102_io_in_b = io_in_b_102; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_103_clock = clock;
  assign FP_multiplier_10ccs_103_reset = reset;
  assign FP_multiplier_10ccs_103_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_103_io_in_b = io_in_b_103; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_104_clock = clock;
  assign FP_multiplier_10ccs_104_reset = reset;
  assign FP_multiplier_10ccs_104_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_104_io_in_b = io_in_b_104; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_105_clock = clock;
  assign FP_multiplier_10ccs_105_reset = reset;
  assign FP_multiplier_10ccs_105_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_105_io_in_b = io_in_b_105; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_106_clock = clock;
  assign FP_multiplier_10ccs_106_reset = reset;
  assign FP_multiplier_10ccs_106_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_106_io_in_b = io_in_b_106; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_107_clock = clock;
  assign FP_multiplier_10ccs_107_reset = reset;
  assign FP_multiplier_10ccs_107_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_107_io_in_b = io_in_b_107; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_108_clock = clock;
  assign FP_multiplier_10ccs_108_reset = reset;
  assign FP_multiplier_10ccs_108_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_108_io_in_b = io_in_b_108; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_109_clock = clock;
  assign FP_multiplier_10ccs_109_reset = reset;
  assign FP_multiplier_10ccs_109_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_109_io_in_b = io_in_b_109; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_110_clock = clock;
  assign FP_multiplier_10ccs_110_reset = reset;
  assign FP_multiplier_10ccs_110_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_110_io_in_b = io_in_b_110; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_111_clock = clock;
  assign FP_multiplier_10ccs_111_reset = reset;
  assign FP_multiplier_10ccs_111_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_111_io_in_b = io_in_b_111; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_112_clock = clock;
  assign FP_multiplier_10ccs_112_reset = reset;
  assign FP_multiplier_10ccs_112_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_112_io_in_b = io_in_b_112; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_113_clock = clock;
  assign FP_multiplier_10ccs_113_reset = reset;
  assign FP_multiplier_10ccs_113_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_113_io_in_b = io_in_b_113; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_114_clock = clock;
  assign FP_multiplier_10ccs_114_reset = reset;
  assign FP_multiplier_10ccs_114_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_114_io_in_b = io_in_b_114; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_115_clock = clock;
  assign FP_multiplier_10ccs_115_reset = reset;
  assign FP_multiplier_10ccs_115_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_115_io_in_b = io_in_b_115; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_116_clock = clock;
  assign FP_multiplier_10ccs_116_reset = reset;
  assign FP_multiplier_10ccs_116_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_116_io_in_b = io_in_b_116; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_117_clock = clock;
  assign FP_multiplier_10ccs_117_reset = reset;
  assign FP_multiplier_10ccs_117_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_117_io_in_b = io_in_b_117; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_118_clock = clock;
  assign FP_multiplier_10ccs_118_reset = reset;
  assign FP_multiplier_10ccs_118_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_118_io_in_b = io_in_b_118; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_119_clock = clock;
  assign FP_multiplier_10ccs_119_reset = reset;
  assign FP_multiplier_10ccs_119_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_119_io_in_b = io_in_b_119; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_120_clock = clock;
  assign FP_multiplier_10ccs_120_reset = reset;
  assign FP_multiplier_10ccs_120_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_120_io_in_b = io_in_b_120; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_121_clock = clock;
  assign FP_multiplier_10ccs_121_reset = reset;
  assign FP_multiplier_10ccs_121_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_121_io_in_b = io_in_b_121; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_122_clock = clock;
  assign FP_multiplier_10ccs_122_reset = reset;
  assign FP_multiplier_10ccs_122_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_122_io_in_b = io_in_b_122; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_123_clock = clock;
  assign FP_multiplier_10ccs_123_reset = reset;
  assign FP_multiplier_10ccs_123_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_123_io_in_b = io_in_b_123; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_124_clock = clock;
  assign FP_multiplier_10ccs_124_reset = reset;
  assign FP_multiplier_10ccs_124_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_124_io_in_b = io_in_b_124; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_125_clock = clock;
  assign FP_multiplier_10ccs_125_reset = reset;
  assign FP_multiplier_10ccs_125_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_125_io_in_b = io_in_b_125; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_126_clock = clock;
  assign FP_multiplier_10ccs_126_reset = reset;
  assign FP_multiplier_10ccs_126_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_126_io_in_b = io_in_b_126; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_multiplier_10ccs_127_clock = clock;
  assign FP_multiplier_10ccs_127_reset = reset;
  assign FP_multiplier_10ccs_127_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2494:30]
  assign FP_multiplier_10ccs_127_io_in_b = io_in_b_127; // @[FloatingPointDesigns.scala 2495:30]
  assign FP_adder_13ccs_clock = clock;
  assign FP_adder_13ccs_reset = reset;
  assign FP_adder_13ccs_io_in_a = FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_io_in_b = FPReg_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_1_clock = clock;
  assign FP_adder_13ccs_1_reset = reset;
  assign FP_adder_13ccs_1_io_in_a = FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_1_io_in_b = FPReg_1_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_2_clock = clock;
  assign FP_adder_13ccs_2_reset = reset;
  assign FP_adder_13ccs_2_io_in_a = FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_2_io_in_b = FPReg_2_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_3_clock = clock;
  assign FP_adder_13ccs_3_reset = reset;
  assign FP_adder_13ccs_3_io_in_a = FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_3_io_in_b = FPReg_3_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_4_clock = clock;
  assign FP_adder_13ccs_4_reset = reset;
  assign FP_adder_13ccs_4_io_in_a = FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_4_io_in_b = FPReg_4_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_5_clock = clock;
  assign FP_adder_13ccs_5_reset = reset;
  assign FP_adder_13ccs_5_io_in_a = FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_5_io_in_b = FPReg_5_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_6_clock = clock;
  assign FP_adder_13ccs_6_reset = reset;
  assign FP_adder_13ccs_6_io_in_a = FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_6_io_in_b = FPReg_6_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_7_clock = clock;
  assign FP_adder_13ccs_7_reset = reset;
  assign FP_adder_13ccs_7_io_in_a = FP_multiplier_10ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_7_io_in_b = FPReg_7_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_8_clock = clock;
  assign FP_adder_13ccs_8_reset = reset;
  assign FP_adder_13ccs_8_io_in_a = FP_multiplier_10ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_8_io_in_b = FPReg_8_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_9_clock = clock;
  assign FP_adder_13ccs_9_reset = reset;
  assign FP_adder_13ccs_9_io_in_a = FP_multiplier_10ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_9_io_in_b = FPReg_9_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_10_clock = clock;
  assign FP_adder_13ccs_10_reset = reset;
  assign FP_adder_13ccs_10_io_in_a = FP_multiplier_10ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_10_io_in_b = FPReg_10_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_11_clock = clock;
  assign FP_adder_13ccs_11_reset = reset;
  assign FP_adder_13ccs_11_io_in_a = FP_multiplier_10ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_11_io_in_b = FPReg_11_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_12_clock = clock;
  assign FP_adder_13ccs_12_reset = reset;
  assign FP_adder_13ccs_12_io_in_a = FP_multiplier_10ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_12_io_in_b = FPReg_12_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_13_clock = clock;
  assign FP_adder_13ccs_13_reset = reset;
  assign FP_adder_13ccs_13_io_in_a = FP_multiplier_10ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_13_io_in_b = FPReg_13_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_14_clock = clock;
  assign FP_adder_13ccs_14_reset = reset;
  assign FP_adder_13ccs_14_io_in_a = FP_multiplier_10ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_14_io_in_b = FPReg_14_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_15_clock = clock;
  assign FP_adder_13ccs_15_reset = reset;
  assign FP_adder_13ccs_15_io_in_a = FP_multiplier_10ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_15_io_in_b = FPReg_15_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_16_clock = clock;
  assign FP_adder_13ccs_16_reset = reset;
  assign FP_adder_13ccs_16_io_in_a = FP_multiplier_10ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_16_io_in_b = FPReg_16_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_17_clock = clock;
  assign FP_adder_13ccs_17_reset = reset;
  assign FP_adder_13ccs_17_io_in_a = FP_multiplier_10ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_17_io_in_b = FPReg_17_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_18_clock = clock;
  assign FP_adder_13ccs_18_reset = reset;
  assign FP_adder_13ccs_18_io_in_a = FP_multiplier_10ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_18_io_in_b = FPReg_18_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_19_clock = clock;
  assign FP_adder_13ccs_19_reset = reset;
  assign FP_adder_13ccs_19_io_in_a = FP_multiplier_10ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_19_io_in_b = FPReg_19_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_20_clock = clock;
  assign FP_adder_13ccs_20_reset = reset;
  assign FP_adder_13ccs_20_io_in_a = FP_multiplier_10ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_20_io_in_b = FPReg_20_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_21_clock = clock;
  assign FP_adder_13ccs_21_reset = reset;
  assign FP_adder_13ccs_21_io_in_a = FP_multiplier_10ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_21_io_in_b = FPReg_21_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_22_clock = clock;
  assign FP_adder_13ccs_22_reset = reset;
  assign FP_adder_13ccs_22_io_in_a = FP_multiplier_10ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_22_io_in_b = FPReg_22_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_23_clock = clock;
  assign FP_adder_13ccs_23_reset = reset;
  assign FP_adder_13ccs_23_io_in_a = FP_multiplier_10ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_23_io_in_b = FPReg_23_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_24_clock = clock;
  assign FP_adder_13ccs_24_reset = reset;
  assign FP_adder_13ccs_24_io_in_a = FP_multiplier_10ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_24_io_in_b = FPReg_24_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_25_clock = clock;
  assign FP_adder_13ccs_25_reset = reset;
  assign FP_adder_13ccs_25_io_in_a = FP_multiplier_10ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_25_io_in_b = FPReg_25_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_26_clock = clock;
  assign FP_adder_13ccs_26_reset = reset;
  assign FP_adder_13ccs_26_io_in_a = FP_multiplier_10ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_26_io_in_b = FPReg_26_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_27_clock = clock;
  assign FP_adder_13ccs_27_reset = reset;
  assign FP_adder_13ccs_27_io_in_a = FP_multiplier_10ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_27_io_in_b = FPReg_27_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_28_clock = clock;
  assign FP_adder_13ccs_28_reset = reset;
  assign FP_adder_13ccs_28_io_in_a = FP_multiplier_10ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_28_io_in_b = FPReg_28_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_29_clock = clock;
  assign FP_adder_13ccs_29_reset = reset;
  assign FP_adder_13ccs_29_io_in_a = FP_multiplier_10ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_29_io_in_b = FPReg_29_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_30_clock = clock;
  assign FP_adder_13ccs_30_reset = reset;
  assign FP_adder_13ccs_30_io_in_a = FP_multiplier_10ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_30_io_in_b = FPReg_30_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_31_clock = clock;
  assign FP_adder_13ccs_31_reset = reset;
  assign FP_adder_13ccs_31_io_in_a = FP_multiplier_10ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_31_io_in_b = FPReg_31_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_32_clock = clock;
  assign FP_adder_13ccs_32_reset = reset;
  assign FP_adder_13ccs_32_io_in_a = FP_multiplier_10ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_32_io_in_b = FPReg_32_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_33_clock = clock;
  assign FP_adder_13ccs_33_reset = reset;
  assign FP_adder_13ccs_33_io_in_a = FP_multiplier_10ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_33_io_in_b = FPReg_33_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_34_clock = clock;
  assign FP_adder_13ccs_34_reset = reset;
  assign FP_adder_13ccs_34_io_in_a = FP_multiplier_10ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_34_io_in_b = FPReg_34_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_35_clock = clock;
  assign FP_adder_13ccs_35_reset = reset;
  assign FP_adder_13ccs_35_io_in_a = FP_multiplier_10ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_35_io_in_b = FPReg_35_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_36_clock = clock;
  assign FP_adder_13ccs_36_reset = reset;
  assign FP_adder_13ccs_36_io_in_a = FP_multiplier_10ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_36_io_in_b = FPReg_36_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_37_clock = clock;
  assign FP_adder_13ccs_37_reset = reset;
  assign FP_adder_13ccs_37_io_in_a = FP_multiplier_10ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_37_io_in_b = FPReg_37_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_38_clock = clock;
  assign FP_adder_13ccs_38_reset = reset;
  assign FP_adder_13ccs_38_io_in_a = FP_multiplier_10ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_38_io_in_b = FPReg_38_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_39_clock = clock;
  assign FP_adder_13ccs_39_reset = reset;
  assign FP_adder_13ccs_39_io_in_a = FP_multiplier_10ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_39_io_in_b = FPReg_39_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_40_clock = clock;
  assign FP_adder_13ccs_40_reset = reset;
  assign FP_adder_13ccs_40_io_in_a = FP_multiplier_10ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_40_io_in_b = FPReg_40_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_41_clock = clock;
  assign FP_adder_13ccs_41_reset = reset;
  assign FP_adder_13ccs_41_io_in_a = FP_multiplier_10ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_41_io_in_b = FPReg_41_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_42_clock = clock;
  assign FP_adder_13ccs_42_reset = reset;
  assign FP_adder_13ccs_42_io_in_a = FP_multiplier_10ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_42_io_in_b = FPReg_42_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_43_clock = clock;
  assign FP_adder_13ccs_43_reset = reset;
  assign FP_adder_13ccs_43_io_in_a = FP_multiplier_10ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_43_io_in_b = FPReg_43_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_44_clock = clock;
  assign FP_adder_13ccs_44_reset = reset;
  assign FP_adder_13ccs_44_io_in_a = FP_multiplier_10ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_44_io_in_b = FPReg_44_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_45_clock = clock;
  assign FP_adder_13ccs_45_reset = reset;
  assign FP_adder_13ccs_45_io_in_a = FP_multiplier_10ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_45_io_in_b = FPReg_45_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_46_clock = clock;
  assign FP_adder_13ccs_46_reset = reset;
  assign FP_adder_13ccs_46_io_in_a = FP_multiplier_10ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_46_io_in_b = FPReg_46_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_47_clock = clock;
  assign FP_adder_13ccs_47_reset = reset;
  assign FP_adder_13ccs_47_io_in_a = FP_multiplier_10ccs_47_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_47_io_in_b = FPReg_47_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_48_clock = clock;
  assign FP_adder_13ccs_48_reset = reset;
  assign FP_adder_13ccs_48_io_in_a = FP_multiplier_10ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_48_io_in_b = FPReg_48_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_49_clock = clock;
  assign FP_adder_13ccs_49_reset = reset;
  assign FP_adder_13ccs_49_io_in_a = FP_multiplier_10ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_49_io_in_b = FPReg_49_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_50_clock = clock;
  assign FP_adder_13ccs_50_reset = reset;
  assign FP_adder_13ccs_50_io_in_a = FP_multiplier_10ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_50_io_in_b = FPReg_50_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_51_clock = clock;
  assign FP_adder_13ccs_51_reset = reset;
  assign FP_adder_13ccs_51_io_in_a = FP_multiplier_10ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_51_io_in_b = FPReg_51_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_52_clock = clock;
  assign FP_adder_13ccs_52_reset = reset;
  assign FP_adder_13ccs_52_io_in_a = FP_multiplier_10ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_52_io_in_b = FPReg_52_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_53_clock = clock;
  assign FP_adder_13ccs_53_reset = reset;
  assign FP_adder_13ccs_53_io_in_a = FP_multiplier_10ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_53_io_in_b = FPReg_53_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_54_clock = clock;
  assign FP_adder_13ccs_54_reset = reset;
  assign FP_adder_13ccs_54_io_in_a = FP_multiplier_10ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_54_io_in_b = FPReg_54_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_55_clock = clock;
  assign FP_adder_13ccs_55_reset = reset;
  assign FP_adder_13ccs_55_io_in_a = FP_multiplier_10ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_55_io_in_b = FPReg_55_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_56_clock = clock;
  assign FP_adder_13ccs_56_reset = reset;
  assign FP_adder_13ccs_56_io_in_a = FP_multiplier_10ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_56_io_in_b = FPReg_56_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_57_clock = clock;
  assign FP_adder_13ccs_57_reset = reset;
  assign FP_adder_13ccs_57_io_in_a = FP_multiplier_10ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_57_io_in_b = FPReg_57_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_58_clock = clock;
  assign FP_adder_13ccs_58_reset = reset;
  assign FP_adder_13ccs_58_io_in_a = FP_multiplier_10ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_58_io_in_b = FPReg_58_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_59_clock = clock;
  assign FP_adder_13ccs_59_reset = reset;
  assign FP_adder_13ccs_59_io_in_a = FP_multiplier_10ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_59_io_in_b = FPReg_59_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_60_clock = clock;
  assign FP_adder_13ccs_60_reset = reset;
  assign FP_adder_13ccs_60_io_in_a = FP_multiplier_10ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_60_io_in_b = FPReg_60_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_61_clock = clock;
  assign FP_adder_13ccs_61_reset = reset;
  assign FP_adder_13ccs_61_io_in_a = FP_multiplier_10ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_61_io_in_b = FPReg_61_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_62_clock = clock;
  assign FP_adder_13ccs_62_reset = reset;
  assign FP_adder_13ccs_62_io_in_a = FP_multiplier_10ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_62_io_in_b = FPReg_62_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_63_clock = clock;
  assign FP_adder_13ccs_63_reset = reset;
  assign FP_adder_13ccs_63_io_in_a = FP_multiplier_10ccs_63_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_63_io_in_b = FPReg_63_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_64_clock = clock;
  assign FP_adder_13ccs_64_reset = reset;
  assign FP_adder_13ccs_64_io_in_a = FP_multiplier_10ccs_64_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_64_io_in_b = FPReg_64_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_65_clock = clock;
  assign FP_adder_13ccs_65_reset = reset;
  assign FP_adder_13ccs_65_io_in_a = FP_multiplier_10ccs_65_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_65_io_in_b = FPReg_65_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_66_clock = clock;
  assign FP_adder_13ccs_66_reset = reset;
  assign FP_adder_13ccs_66_io_in_a = FP_multiplier_10ccs_66_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_66_io_in_b = FPReg_66_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_67_clock = clock;
  assign FP_adder_13ccs_67_reset = reset;
  assign FP_adder_13ccs_67_io_in_a = FP_multiplier_10ccs_67_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_67_io_in_b = FPReg_67_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_68_clock = clock;
  assign FP_adder_13ccs_68_reset = reset;
  assign FP_adder_13ccs_68_io_in_a = FP_multiplier_10ccs_68_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_68_io_in_b = FPReg_68_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_69_clock = clock;
  assign FP_adder_13ccs_69_reset = reset;
  assign FP_adder_13ccs_69_io_in_a = FP_multiplier_10ccs_69_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_69_io_in_b = FPReg_69_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_70_clock = clock;
  assign FP_adder_13ccs_70_reset = reset;
  assign FP_adder_13ccs_70_io_in_a = FP_multiplier_10ccs_70_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_70_io_in_b = FPReg_70_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_71_clock = clock;
  assign FP_adder_13ccs_71_reset = reset;
  assign FP_adder_13ccs_71_io_in_a = FP_multiplier_10ccs_71_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_71_io_in_b = FPReg_71_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_72_clock = clock;
  assign FP_adder_13ccs_72_reset = reset;
  assign FP_adder_13ccs_72_io_in_a = FP_multiplier_10ccs_72_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_72_io_in_b = FPReg_72_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_73_clock = clock;
  assign FP_adder_13ccs_73_reset = reset;
  assign FP_adder_13ccs_73_io_in_a = FP_multiplier_10ccs_73_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_73_io_in_b = FPReg_73_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_74_clock = clock;
  assign FP_adder_13ccs_74_reset = reset;
  assign FP_adder_13ccs_74_io_in_a = FP_multiplier_10ccs_74_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_74_io_in_b = FPReg_74_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_75_clock = clock;
  assign FP_adder_13ccs_75_reset = reset;
  assign FP_adder_13ccs_75_io_in_a = FP_multiplier_10ccs_75_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_75_io_in_b = FPReg_75_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_76_clock = clock;
  assign FP_adder_13ccs_76_reset = reset;
  assign FP_adder_13ccs_76_io_in_a = FP_multiplier_10ccs_76_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_76_io_in_b = FPReg_76_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_77_clock = clock;
  assign FP_adder_13ccs_77_reset = reset;
  assign FP_adder_13ccs_77_io_in_a = FP_multiplier_10ccs_77_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_77_io_in_b = FPReg_77_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_78_clock = clock;
  assign FP_adder_13ccs_78_reset = reset;
  assign FP_adder_13ccs_78_io_in_a = FP_multiplier_10ccs_78_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_78_io_in_b = FPReg_78_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_79_clock = clock;
  assign FP_adder_13ccs_79_reset = reset;
  assign FP_adder_13ccs_79_io_in_a = FP_multiplier_10ccs_79_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_79_io_in_b = FPReg_79_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_80_clock = clock;
  assign FP_adder_13ccs_80_reset = reset;
  assign FP_adder_13ccs_80_io_in_a = FP_multiplier_10ccs_80_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_80_io_in_b = FPReg_80_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_81_clock = clock;
  assign FP_adder_13ccs_81_reset = reset;
  assign FP_adder_13ccs_81_io_in_a = FP_multiplier_10ccs_81_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_81_io_in_b = FPReg_81_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_82_clock = clock;
  assign FP_adder_13ccs_82_reset = reset;
  assign FP_adder_13ccs_82_io_in_a = FP_multiplier_10ccs_82_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_82_io_in_b = FPReg_82_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_83_clock = clock;
  assign FP_adder_13ccs_83_reset = reset;
  assign FP_adder_13ccs_83_io_in_a = FP_multiplier_10ccs_83_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_83_io_in_b = FPReg_83_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_84_clock = clock;
  assign FP_adder_13ccs_84_reset = reset;
  assign FP_adder_13ccs_84_io_in_a = FP_multiplier_10ccs_84_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_84_io_in_b = FPReg_84_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_85_clock = clock;
  assign FP_adder_13ccs_85_reset = reset;
  assign FP_adder_13ccs_85_io_in_a = FP_multiplier_10ccs_85_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_85_io_in_b = FPReg_85_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_86_clock = clock;
  assign FP_adder_13ccs_86_reset = reset;
  assign FP_adder_13ccs_86_io_in_a = FP_multiplier_10ccs_86_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_86_io_in_b = FPReg_86_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_87_clock = clock;
  assign FP_adder_13ccs_87_reset = reset;
  assign FP_adder_13ccs_87_io_in_a = FP_multiplier_10ccs_87_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_87_io_in_b = FPReg_87_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_88_clock = clock;
  assign FP_adder_13ccs_88_reset = reset;
  assign FP_adder_13ccs_88_io_in_a = FP_multiplier_10ccs_88_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_88_io_in_b = FPReg_88_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_89_clock = clock;
  assign FP_adder_13ccs_89_reset = reset;
  assign FP_adder_13ccs_89_io_in_a = FP_multiplier_10ccs_89_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_89_io_in_b = FPReg_89_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_90_clock = clock;
  assign FP_adder_13ccs_90_reset = reset;
  assign FP_adder_13ccs_90_io_in_a = FP_multiplier_10ccs_90_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_90_io_in_b = FPReg_90_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_91_clock = clock;
  assign FP_adder_13ccs_91_reset = reset;
  assign FP_adder_13ccs_91_io_in_a = FP_multiplier_10ccs_91_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_91_io_in_b = FPReg_91_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_92_clock = clock;
  assign FP_adder_13ccs_92_reset = reset;
  assign FP_adder_13ccs_92_io_in_a = FP_multiplier_10ccs_92_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_92_io_in_b = FPReg_92_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_93_clock = clock;
  assign FP_adder_13ccs_93_reset = reset;
  assign FP_adder_13ccs_93_io_in_a = FP_multiplier_10ccs_93_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_93_io_in_b = FPReg_93_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_94_clock = clock;
  assign FP_adder_13ccs_94_reset = reset;
  assign FP_adder_13ccs_94_io_in_a = FP_multiplier_10ccs_94_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_94_io_in_b = FPReg_94_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_95_clock = clock;
  assign FP_adder_13ccs_95_reset = reset;
  assign FP_adder_13ccs_95_io_in_a = FP_multiplier_10ccs_95_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_95_io_in_b = FPReg_95_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_96_clock = clock;
  assign FP_adder_13ccs_96_reset = reset;
  assign FP_adder_13ccs_96_io_in_a = FP_multiplier_10ccs_96_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_96_io_in_b = FPReg_96_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_97_clock = clock;
  assign FP_adder_13ccs_97_reset = reset;
  assign FP_adder_13ccs_97_io_in_a = FP_multiplier_10ccs_97_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_97_io_in_b = FPReg_97_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_98_clock = clock;
  assign FP_adder_13ccs_98_reset = reset;
  assign FP_adder_13ccs_98_io_in_a = FP_multiplier_10ccs_98_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_98_io_in_b = FPReg_98_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_99_clock = clock;
  assign FP_adder_13ccs_99_reset = reset;
  assign FP_adder_13ccs_99_io_in_a = FP_multiplier_10ccs_99_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_99_io_in_b = FPReg_99_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_100_clock = clock;
  assign FP_adder_13ccs_100_reset = reset;
  assign FP_adder_13ccs_100_io_in_a = FP_multiplier_10ccs_100_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_100_io_in_b = FPReg_100_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_101_clock = clock;
  assign FP_adder_13ccs_101_reset = reset;
  assign FP_adder_13ccs_101_io_in_a = FP_multiplier_10ccs_101_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_101_io_in_b = FPReg_101_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_102_clock = clock;
  assign FP_adder_13ccs_102_reset = reset;
  assign FP_adder_13ccs_102_io_in_a = FP_multiplier_10ccs_102_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_102_io_in_b = FPReg_102_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_103_clock = clock;
  assign FP_adder_13ccs_103_reset = reset;
  assign FP_adder_13ccs_103_io_in_a = FP_multiplier_10ccs_103_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_103_io_in_b = FPReg_103_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_104_clock = clock;
  assign FP_adder_13ccs_104_reset = reset;
  assign FP_adder_13ccs_104_io_in_a = FP_multiplier_10ccs_104_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_104_io_in_b = FPReg_104_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_105_clock = clock;
  assign FP_adder_13ccs_105_reset = reset;
  assign FP_adder_13ccs_105_io_in_a = FP_multiplier_10ccs_105_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_105_io_in_b = FPReg_105_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_106_clock = clock;
  assign FP_adder_13ccs_106_reset = reset;
  assign FP_adder_13ccs_106_io_in_a = FP_multiplier_10ccs_106_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_106_io_in_b = FPReg_106_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_107_clock = clock;
  assign FP_adder_13ccs_107_reset = reset;
  assign FP_adder_13ccs_107_io_in_a = FP_multiplier_10ccs_107_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_107_io_in_b = FPReg_107_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_108_clock = clock;
  assign FP_adder_13ccs_108_reset = reset;
  assign FP_adder_13ccs_108_io_in_a = FP_multiplier_10ccs_108_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_108_io_in_b = FPReg_108_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_109_clock = clock;
  assign FP_adder_13ccs_109_reset = reset;
  assign FP_adder_13ccs_109_io_in_a = FP_multiplier_10ccs_109_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_109_io_in_b = FPReg_109_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_110_clock = clock;
  assign FP_adder_13ccs_110_reset = reset;
  assign FP_adder_13ccs_110_io_in_a = FP_multiplier_10ccs_110_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_110_io_in_b = FPReg_110_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_111_clock = clock;
  assign FP_adder_13ccs_111_reset = reset;
  assign FP_adder_13ccs_111_io_in_a = FP_multiplier_10ccs_111_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_111_io_in_b = FPReg_111_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_112_clock = clock;
  assign FP_adder_13ccs_112_reset = reset;
  assign FP_adder_13ccs_112_io_in_a = FP_multiplier_10ccs_112_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_112_io_in_b = FPReg_112_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_113_clock = clock;
  assign FP_adder_13ccs_113_reset = reset;
  assign FP_adder_13ccs_113_io_in_a = FP_multiplier_10ccs_113_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_113_io_in_b = FPReg_113_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_114_clock = clock;
  assign FP_adder_13ccs_114_reset = reset;
  assign FP_adder_13ccs_114_io_in_a = FP_multiplier_10ccs_114_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_114_io_in_b = FPReg_114_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_115_clock = clock;
  assign FP_adder_13ccs_115_reset = reset;
  assign FP_adder_13ccs_115_io_in_a = FP_multiplier_10ccs_115_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_115_io_in_b = FPReg_115_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_116_clock = clock;
  assign FP_adder_13ccs_116_reset = reset;
  assign FP_adder_13ccs_116_io_in_a = FP_multiplier_10ccs_116_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_116_io_in_b = FPReg_116_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_117_clock = clock;
  assign FP_adder_13ccs_117_reset = reset;
  assign FP_adder_13ccs_117_io_in_a = FP_multiplier_10ccs_117_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_117_io_in_b = FPReg_117_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_118_clock = clock;
  assign FP_adder_13ccs_118_reset = reset;
  assign FP_adder_13ccs_118_io_in_a = FP_multiplier_10ccs_118_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_118_io_in_b = FPReg_118_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_119_clock = clock;
  assign FP_adder_13ccs_119_reset = reset;
  assign FP_adder_13ccs_119_io_in_a = FP_multiplier_10ccs_119_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_119_io_in_b = FPReg_119_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_120_clock = clock;
  assign FP_adder_13ccs_120_reset = reset;
  assign FP_adder_13ccs_120_io_in_a = FP_multiplier_10ccs_120_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_120_io_in_b = FPReg_120_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_121_clock = clock;
  assign FP_adder_13ccs_121_reset = reset;
  assign FP_adder_13ccs_121_io_in_a = FP_multiplier_10ccs_121_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_121_io_in_b = FPReg_121_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_122_clock = clock;
  assign FP_adder_13ccs_122_reset = reset;
  assign FP_adder_13ccs_122_io_in_a = FP_multiplier_10ccs_122_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_122_io_in_b = FPReg_122_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_123_clock = clock;
  assign FP_adder_13ccs_123_reset = reset;
  assign FP_adder_13ccs_123_io_in_a = FP_multiplier_10ccs_123_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_123_io_in_b = FPReg_123_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_124_clock = clock;
  assign FP_adder_13ccs_124_reset = reset;
  assign FP_adder_13ccs_124_io_in_a = FP_multiplier_10ccs_124_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_124_io_in_b = FPReg_124_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_125_clock = clock;
  assign FP_adder_13ccs_125_reset = reset;
  assign FP_adder_13ccs_125_io_in_a = FP_multiplier_10ccs_125_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_125_io_in_b = FPReg_125_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_126_clock = clock;
  assign FP_adder_13ccs_126_reset = reset;
  assign FP_adder_13ccs_126_io_in_a = FP_multiplier_10ccs_126_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_126_io_in_b = FPReg_126_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FP_adder_13ccs_127_clock = clock;
  assign FP_adder_13ccs_127_reset = reset;
  assign FP_adder_13ccs_127_io_in_a = FP_multiplier_10ccs_127_io_out_s; // @[FloatingPointDesigns.scala 2497:27]
  assign FP_adder_13ccs_127_io_in_b = FPReg_127_io_out; // @[FloatingPointDesigns.scala 2498:27]
  assign FPReg_clock = clock;
  assign FPReg_reset = reset;
  assign FPReg_io_in = io_in_c_0; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_1_clock = clock;
  assign FPReg_1_reset = reset;
  assign FPReg_1_io_in = io_in_c_1; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_2_clock = clock;
  assign FPReg_2_reset = reset;
  assign FPReg_2_io_in = io_in_c_2; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_3_clock = clock;
  assign FPReg_3_reset = reset;
  assign FPReg_3_io_in = io_in_c_3; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_4_clock = clock;
  assign FPReg_4_reset = reset;
  assign FPReg_4_io_in = io_in_c_4; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_5_clock = clock;
  assign FPReg_5_reset = reset;
  assign FPReg_5_io_in = io_in_c_5; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_6_clock = clock;
  assign FPReg_6_reset = reset;
  assign FPReg_6_io_in = io_in_c_6; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_7_clock = clock;
  assign FPReg_7_reset = reset;
  assign FPReg_7_io_in = io_in_c_7; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_8_clock = clock;
  assign FPReg_8_reset = reset;
  assign FPReg_8_io_in = io_in_c_8; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_9_clock = clock;
  assign FPReg_9_reset = reset;
  assign FPReg_9_io_in = io_in_c_9; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_10_clock = clock;
  assign FPReg_10_reset = reset;
  assign FPReg_10_io_in = io_in_c_10; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_11_clock = clock;
  assign FPReg_11_reset = reset;
  assign FPReg_11_io_in = io_in_c_11; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_12_clock = clock;
  assign FPReg_12_reset = reset;
  assign FPReg_12_io_in = io_in_c_12; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_13_clock = clock;
  assign FPReg_13_reset = reset;
  assign FPReg_13_io_in = io_in_c_13; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_14_clock = clock;
  assign FPReg_14_reset = reset;
  assign FPReg_14_io_in = io_in_c_14; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_15_clock = clock;
  assign FPReg_15_reset = reset;
  assign FPReg_15_io_in = io_in_c_15; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_16_clock = clock;
  assign FPReg_16_reset = reset;
  assign FPReg_16_io_in = io_in_c_16; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_17_clock = clock;
  assign FPReg_17_reset = reset;
  assign FPReg_17_io_in = io_in_c_17; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_18_clock = clock;
  assign FPReg_18_reset = reset;
  assign FPReg_18_io_in = io_in_c_18; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_19_clock = clock;
  assign FPReg_19_reset = reset;
  assign FPReg_19_io_in = io_in_c_19; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_20_clock = clock;
  assign FPReg_20_reset = reset;
  assign FPReg_20_io_in = io_in_c_20; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_21_clock = clock;
  assign FPReg_21_reset = reset;
  assign FPReg_21_io_in = io_in_c_21; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_22_clock = clock;
  assign FPReg_22_reset = reset;
  assign FPReg_22_io_in = io_in_c_22; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_23_clock = clock;
  assign FPReg_23_reset = reset;
  assign FPReg_23_io_in = io_in_c_23; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_24_clock = clock;
  assign FPReg_24_reset = reset;
  assign FPReg_24_io_in = io_in_c_24; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_25_clock = clock;
  assign FPReg_25_reset = reset;
  assign FPReg_25_io_in = io_in_c_25; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_26_clock = clock;
  assign FPReg_26_reset = reset;
  assign FPReg_26_io_in = io_in_c_26; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_27_clock = clock;
  assign FPReg_27_reset = reset;
  assign FPReg_27_io_in = io_in_c_27; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_28_clock = clock;
  assign FPReg_28_reset = reset;
  assign FPReg_28_io_in = io_in_c_28; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_29_clock = clock;
  assign FPReg_29_reset = reset;
  assign FPReg_29_io_in = io_in_c_29; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_30_clock = clock;
  assign FPReg_30_reset = reset;
  assign FPReg_30_io_in = io_in_c_30; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_31_clock = clock;
  assign FPReg_31_reset = reset;
  assign FPReg_31_io_in = io_in_c_31; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_32_clock = clock;
  assign FPReg_32_reset = reset;
  assign FPReg_32_io_in = io_in_c_32; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_33_clock = clock;
  assign FPReg_33_reset = reset;
  assign FPReg_33_io_in = io_in_c_33; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_34_clock = clock;
  assign FPReg_34_reset = reset;
  assign FPReg_34_io_in = io_in_c_34; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_35_clock = clock;
  assign FPReg_35_reset = reset;
  assign FPReg_35_io_in = io_in_c_35; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_36_clock = clock;
  assign FPReg_36_reset = reset;
  assign FPReg_36_io_in = io_in_c_36; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_37_clock = clock;
  assign FPReg_37_reset = reset;
  assign FPReg_37_io_in = io_in_c_37; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_38_clock = clock;
  assign FPReg_38_reset = reset;
  assign FPReg_38_io_in = io_in_c_38; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_39_clock = clock;
  assign FPReg_39_reset = reset;
  assign FPReg_39_io_in = io_in_c_39; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_40_clock = clock;
  assign FPReg_40_reset = reset;
  assign FPReg_40_io_in = io_in_c_40; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_41_clock = clock;
  assign FPReg_41_reset = reset;
  assign FPReg_41_io_in = io_in_c_41; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_42_clock = clock;
  assign FPReg_42_reset = reset;
  assign FPReg_42_io_in = io_in_c_42; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_43_clock = clock;
  assign FPReg_43_reset = reset;
  assign FPReg_43_io_in = io_in_c_43; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_44_clock = clock;
  assign FPReg_44_reset = reset;
  assign FPReg_44_io_in = io_in_c_44; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_45_clock = clock;
  assign FPReg_45_reset = reset;
  assign FPReg_45_io_in = io_in_c_45; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_46_clock = clock;
  assign FPReg_46_reset = reset;
  assign FPReg_46_io_in = io_in_c_46; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_47_clock = clock;
  assign FPReg_47_reset = reset;
  assign FPReg_47_io_in = io_in_c_47; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_48_clock = clock;
  assign FPReg_48_reset = reset;
  assign FPReg_48_io_in = io_in_c_48; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_49_clock = clock;
  assign FPReg_49_reset = reset;
  assign FPReg_49_io_in = io_in_c_49; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_50_clock = clock;
  assign FPReg_50_reset = reset;
  assign FPReg_50_io_in = io_in_c_50; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_51_clock = clock;
  assign FPReg_51_reset = reset;
  assign FPReg_51_io_in = io_in_c_51; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_52_clock = clock;
  assign FPReg_52_reset = reset;
  assign FPReg_52_io_in = io_in_c_52; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_53_clock = clock;
  assign FPReg_53_reset = reset;
  assign FPReg_53_io_in = io_in_c_53; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_54_clock = clock;
  assign FPReg_54_reset = reset;
  assign FPReg_54_io_in = io_in_c_54; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_55_clock = clock;
  assign FPReg_55_reset = reset;
  assign FPReg_55_io_in = io_in_c_55; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_56_clock = clock;
  assign FPReg_56_reset = reset;
  assign FPReg_56_io_in = io_in_c_56; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_57_clock = clock;
  assign FPReg_57_reset = reset;
  assign FPReg_57_io_in = io_in_c_57; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_58_clock = clock;
  assign FPReg_58_reset = reset;
  assign FPReg_58_io_in = io_in_c_58; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_59_clock = clock;
  assign FPReg_59_reset = reset;
  assign FPReg_59_io_in = io_in_c_59; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_60_clock = clock;
  assign FPReg_60_reset = reset;
  assign FPReg_60_io_in = io_in_c_60; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_61_clock = clock;
  assign FPReg_61_reset = reset;
  assign FPReg_61_io_in = io_in_c_61; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_62_clock = clock;
  assign FPReg_62_reset = reset;
  assign FPReg_62_io_in = io_in_c_62; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_63_clock = clock;
  assign FPReg_63_reset = reset;
  assign FPReg_63_io_in = io_in_c_63; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_64_clock = clock;
  assign FPReg_64_reset = reset;
  assign FPReg_64_io_in = io_in_c_64; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_65_clock = clock;
  assign FPReg_65_reset = reset;
  assign FPReg_65_io_in = io_in_c_65; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_66_clock = clock;
  assign FPReg_66_reset = reset;
  assign FPReg_66_io_in = io_in_c_66; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_67_clock = clock;
  assign FPReg_67_reset = reset;
  assign FPReg_67_io_in = io_in_c_67; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_68_clock = clock;
  assign FPReg_68_reset = reset;
  assign FPReg_68_io_in = io_in_c_68; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_69_clock = clock;
  assign FPReg_69_reset = reset;
  assign FPReg_69_io_in = io_in_c_69; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_70_clock = clock;
  assign FPReg_70_reset = reset;
  assign FPReg_70_io_in = io_in_c_70; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_71_clock = clock;
  assign FPReg_71_reset = reset;
  assign FPReg_71_io_in = io_in_c_71; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_72_clock = clock;
  assign FPReg_72_reset = reset;
  assign FPReg_72_io_in = io_in_c_72; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_73_clock = clock;
  assign FPReg_73_reset = reset;
  assign FPReg_73_io_in = io_in_c_73; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_74_clock = clock;
  assign FPReg_74_reset = reset;
  assign FPReg_74_io_in = io_in_c_74; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_75_clock = clock;
  assign FPReg_75_reset = reset;
  assign FPReg_75_io_in = io_in_c_75; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_76_clock = clock;
  assign FPReg_76_reset = reset;
  assign FPReg_76_io_in = io_in_c_76; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_77_clock = clock;
  assign FPReg_77_reset = reset;
  assign FPReg_77_io_in = io_in_c_77; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_78_clock = clock;
  assign FPReg_78_reset = reset;
  assign FPReg_78_io_in = io_in_c_78; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_79_clock = clock;
  assign FPReg_79_reset = reset;
  assign FPReg_79_io_in = io_in_c_79; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_80_clock = clock;
  assign FPReg_80_reset = reset;
  assign FPReg_80_io_in = io_in_c_80; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_81_clock = clock;
  assign FPReg_81_reset = reset;
  assign FPReg_81_io_in = io_in_c_81; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_82_clock = clock;
  assign FPReg_82_reset = reset;
  assign FPReg_82_io_in = io_in_c_82; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_83_clock = clock;
  assign FPReg_83_reset = reset;
  assign FPReg_83_io_in = io_in_c_83; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_84_clock = clock;
  assign FPReg_84_reset = reset;
  assign FPReg_84_io_in = io_in_c_84; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_85_clock = clock;
  assign FPReg_85_reset = reset;
  assign FPReg_85_io_in = io_in_c_85; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_86_clock = clock;
  assign FPReg_86_reset = reset;
  assign FPReg_86_io_in = io_in_c_86; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_87_clock = clock;
  assign FPReg_87_reset = reset;
  assign FPReg_87_io_in = io_in_c_87; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_88_clock = clock;
  assign FPReg_88_reset = reset;
  assign FPReg_88_io_in = io_in_c_88; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_89_clock = clock;
  assign FPReg_89_reset = reset;
  assign FPReg_89_io_in = io_in_c_89; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_90_clock = clock;
  assign FPReg_90_reset = reset;
  assign FPReg_90_io_in = io_in_c_90; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_91_clock = clock;
  assign FPReg_91_reset = reset;
  assign FPReg_91_io_in = io_in_c_91; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_92_clock = clock;
  assign FPReg_92_reset = reset;
  assign FPReg_92_io_in = io_in_c_92; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_93_clock = clock;
  assign FPReg_93_reset = reset;
  assign FPReg_93_io_in = io_in_c_93; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_94_clock = clock;
  assign FPReg_94_reset = reset;
  assign FPReg_94_io_in = io_in_c_94; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_95_clock = clock;
  assign FPReg_95_reset = reset;
  assign FPReg_95_io_in = io_in_c_95; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_96_clock = clock;
  assign FPReg_96_reset = reset;
  assign FPReg_96_io_in = io_in_c_96; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_97_clock = clock;
  assign FPReg_97_reset = reset;
  assign FPReg_97_io_in = io_in_c_97; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_98_clock = clock;
  assign FPReg_98_reset = reset;
  assign FPReg_98_io_in = io_in_c_98; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_99_clock = clock;
  assign FPReg_99_reset = reset;
  assign FPReg_99_io_in = io_in_c_99; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_100_clock = clock;
  assign FPReg_100_reset = reset;
  assign FPReg_100_io_in = io_in_c_100; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_101_clock = clock;
  assign FPReg_101_reset = reset;
  assign FPReg_101_io_in = io_in_c_101; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_102_clock = clock;
  assign FPReg_102_reset = reset;
  assign FPReg_102_io_in = io_in_c_102; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_103_clock = clock;
  assign FPReg_103_reset = reset;
  assign FPReg_103_io_in = io_in_c_103; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_104_clock = clock;
  assign FPReg_104_reset = reset;
  assign FPReg_104_io_in = io_in_c_104; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_105_clock = clock;
  assign FPReg_105_reset = reset;
  assign FPReg_105_io_in = io_in_c_105; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_106_clock = clock;
  assign FPReg_106_reset = reset;
  assign FPReg_106_io_in = io_in_c_106; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_107_clock = clock;
  assign FPReg_107_reset = reset;
  assign FPReg_107_io_in = io_in_c_107; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_108_clock = clock;
  assign FPReg_108_reset = reset;
  assign FPReg_108_io_in = io_in_c_108; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_109_clock = clock;
  assign FPReg_109_reset = reset;
  assign FPReg_109_io_in = io_in_c_109; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_110_clock = clock;
  assign FPReg_110_reset = reset;
  assign FPReg_110_io_in = io_in_c_110; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_111_clock = clock;
  assign FPReg_111_reset = reset;
  assign FPReg_111_io_in = io_in_c_111; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_112_clock = clock;
  assign FPReg_112_reset = reset;
  assign FPReg_112_io_in = io_in_c_112; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_113_clock = clock;
  assign FPReg_113_reset = reset;
  assign FPReg_113_io_in = io_in_c_113; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_114_clock = clock;
  assign FPReg_114_reset = reset;
  assign FPReg_114_io_in = io_in_c_114; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_115_clock = clock;
  assign FPReg_115_reset = reset;
  assign FPReg_115_io_in = io_in_c_115; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_116_clock = clock;
  assign FPReg_116_reset = reset;
  assign FPReg_116_io_in = io_in_c_116; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_117_clock = clock;
  assign FPReg_117_reset = reset;
  assign FPReg_117_io_in = io_in_c_117; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_118_clock = clock;
  assign FPReg_118_reset = reset;
  assign FPReg_118_io_in = io_in_c_118; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_119_clock = clock;
  assign FPReg_119_reset = reset;
  assign FPReg_119_io_in = io_in_c_119; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_120_clock = clock;
  assign FPReg_120_reset = reset;
  assign FPReg_120_io_in = io_in_c_120; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_121_clock = clock;
  assign FPReg_121_reset = reset;
  assign FPReg_121_io_in = io_in_c_121; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_122_clock = clock;
  assign FPReg_122_reset = reset;
  assign FPReg_122_io_in = io_in_c_122; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_123_clock = clock;
  assign FPReg_123_reset = reset;
  assign FPReg_123_io_in = io_in_c_123; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_124_clock = clock;
  assign FPReg_124_reset = reset;
  assign FPReg_124_io_in = io_in_c_124; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_125_clock = clock;
  assign FPReg_125_reset = reset;
  assign FPReg_125_io_in = io_in_c_125; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_126_clock = clock;
  assign FPReg_126_reset = reset;
  assign FPReg_126_io_in = io_in_c_126; // @[FloatingPointDesigns.scala 2496:25]
  assign FPReg_127_clock = clock;
  assign FPReg_127_reset = reset;
  assign FPReg_127_io_in = io_in_c_127; // @[FloatingPointDesigns.scala 2496:25]
endmodule
module hh_datapath_1(
  input           io_clk,
  input           io_rst,
  input  [15:0]   io_hh_cnt,
  input           io_d1_rdy,
  input           io_d1_vld,
  input           io_d2_vld,
  input           io_vk1_vld,
  input           io_d3_rdy,
  input           io_d3_vld,
  input           io_tk_vld,
  input           io_d4_rdy,
  input           io_d5_rdy,
  input           io_d5_vld,
  input           io_yj_sft,
  input           io_d4_sft,
  input  [4095:0] io_hh_din,
  output [4095:0] io_hh_dout
);
`ifdef RANDOMIZE_REG_INIT
  reg [4095:0] _RAND_0;
  reg [243711:0] _RAND_1;
  reg [243711:0] _RAND_2;
  reg [243711:0] _RAND_3;
  reg [243711:0] _RAND_4;
  reg [4095:0] _RAND_5;
  reg [4095:0] _RAND_6;
  reg [4095:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [4063:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  FP_DDOT_dp_clock; // @[hh_datapath_chisel.scala 248:21]
  wire  FP_DDOT_dp_reset; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_0; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_1; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_2; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_3; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_4; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_5; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_6; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_7; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_8; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_9; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_10; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_11; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_12; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_13; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_14; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_15; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_16; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_17; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_18; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_19; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_20; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_21; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_22; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_23; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_24; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_25; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_26; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_27; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_28; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_29; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_30; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_31; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_32; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_33; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_34; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_35; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_36; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_37; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_38; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_39; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_40; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_41; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_42; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_43; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_44; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_45; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_46; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_47; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_48; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_49; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_50; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_51; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_52; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_53; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_54; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_55; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_56; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_57; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_58; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_59; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_60; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_61; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_62; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_63; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_64; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_65; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_66; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_67; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_68; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_69; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_70; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_71; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_72; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_73; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_74; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_75; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_76; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_77; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_78; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_79; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_80; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_81; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_82; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_83; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_84; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_85; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_86; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_87; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_88; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_89; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_90; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_91; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_92; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_93; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_94; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_95; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_96; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_97; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_98; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_99; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_100; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_101; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_102; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_103; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_104; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_105; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_106; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_107; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_108; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_109; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_110; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_111; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_112; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_113; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_114; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_115; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_116; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_117; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_118; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_119; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_120; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_121; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_122; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_123; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_124; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_125; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_126; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_127; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_0; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_1; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_2; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_3; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_4; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_5; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_6; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_7; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_8; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_9; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_10; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_11; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_12; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_13; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_14; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_15; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_16; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_17; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_18; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_19; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_20; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_21; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_22; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_23; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_24; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_25; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_26; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_27; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_28; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_29; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_30; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_31; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_32; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_33; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_34; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_35; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_36; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_37; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_38; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_39; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_40; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_41; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_42; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_43; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_44; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_45; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_46; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_47; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_48; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_49; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_50; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_51; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_52; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_53; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_54; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_55; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_56; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_57; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_58; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_59; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_60; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_61; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_62; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_63; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_64; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_65; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_66; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_67; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_68; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_69; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_70; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_71; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_72; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_73; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_74; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_75; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_76; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_77; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_78; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_79; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_80; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_81; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_82; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_83; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_84; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_85; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_86; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_87; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_88; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_89; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_90; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_91; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_92; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_93; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_94; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_95; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_96; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_97; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_98; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_99; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_100; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_101; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_102; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_103; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_104; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_105; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_106; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_107; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_108; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_109; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_110; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_111; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_112; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_113; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_114; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_115; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_116; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_117; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_118; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_119; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_120; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_121; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_122; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_123; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_124; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_125; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_126; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_127; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_out_s; // @[hh_datapath_chisel.scala 248:21]
  wire  FP_square_root_newfpu_clock; // @[hh_datapath_chisel.scala 256:22]
  wire  FP_square_root_newfpu_reset; // @[hh_datapath_chisel.scala 256:22]
  wire [31:0] FP_square_root_newfpu_io_in_a; // @[hh_datapath_chisel.scala 256:22]
  wire [31:0] FP_square_root_newfpu_io_out_s; // @[hh_datapath_chisel.scala 256:22]
  wire  hqr5_clock; // @[hh_datapath_chisel.scala 261:20]
  wire  hqr5_reset; // @[hh_datapath_chisel.scala 261:20]
  wire [31:0] hqr5_io_in_a; // @[hh_datapath_chisel.scala 261:20]
  wire [31:0] hqr5_io_in_b; // @[hh_datapath_chisel.scala 261:20]
  wire [31:0] hqr5_io_out_s; // @[hh_datapath_chisel.scala 261:20]
  wire  hqr7_clock; // @[hh_datapath_chisel.scala 266:20]
  wire  hqr7_reset; // @[hh_datapath_chisel.scala 266:20]
  wire [31:0] hqr7_io_in_a; // @[hh_datapath_chisel.scala 266:20]
  wire [31:0] hqr7_io_out_s; // @[hh_datapath_chisel.scala 266:20]
  wire  FP_multiplier_10ccs_clock; // @[hh_datapath_chisel.scala 270:21]
  wire  FP_multiplier_10ccs_reset; // @[hh_datapath_chisel.scala 270:21]
  wire [31:0] FP_multiplier_10ccs_io_in_a; // @[hh_datapath_chisel.scala 270:21]
  wire [31:0] FP_multiplier_10ccs_io_in_b; // @[hh_datapath_chisel.scala 270:21]
  wire [31:0] FP_multiplier_10ccs_io_out_s; // @[hh_datapath_chisel.scala 270:21]
  wire  axpy_dp_clock; // @[hh_datapath_chisel.scala 276:20]
  wire  axpy_dp_reset; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_a; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_0; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_1; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_2; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_3; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_4; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_5; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_6; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_7; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_8; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_9; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_10; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_11; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_12; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_13; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_14; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_15; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_16; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_17; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_18; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_19; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_20; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_21; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_22; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_23; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_24; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_25; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_26; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_27; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_28; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_29; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_30; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_31; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_32; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_33; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_34; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_35; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_36; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_37; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_38; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_39; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_40; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_41; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_42; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_43; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_44; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_45; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_46; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_47; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_48; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_49; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_50; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_51; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_52; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_53; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_54; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_55; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_56; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_57; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_58; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_59; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_60; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_61; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_62; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_63; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_64; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_65; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_66; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_67; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_68; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_69; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_70; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_71; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_72; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_73; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_74; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_75; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_76; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_77; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_78; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_79; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_80; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_81; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_82; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_83; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_84; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_85; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_86; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_87; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_88; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_89; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_90; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_91; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_92; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_93; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_94; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_95; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_96; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_97; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_98; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_99; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_100; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_101; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_102; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_103; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_104; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_105; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_106; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_107; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_108; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_109; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_110; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_111; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_112; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_113; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_114; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_115; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_116; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_117; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_118; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_119; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_120; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_121; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_122; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_123; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_124; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_125; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_126; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_127; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_0; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_1; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_2; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_3; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_4; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_5; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_6; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_7; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_8; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_9; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_10; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_11; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_12; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_13; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_14; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_15; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_16; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_17; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_18; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_19; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_20; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_21; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_22; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_23; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_24; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_25; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_26; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_27; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_28; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_29; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_30; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_31; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_32; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_33; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_34; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_35; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_36; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_37; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_38; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_39; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_40; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_41; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_42; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_43; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_44; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_45; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_46; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_47; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_48; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_49; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_50; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_51; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_52; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_53; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_54; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_55; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_56; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_57; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_58; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_59; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_60; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_61; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_62; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_63; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_64; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_65; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_66; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_67; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_68; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_69; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_70; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_71; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_72; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_73; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_74; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_75; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_76; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_77; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_78; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_79; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_80; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_81; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_82; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_83; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_84; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_85; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_86; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_87; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_88; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_89; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_90; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_91; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_92; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_93; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_94; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_95; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_96; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_97; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_98; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_99; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_100; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_101; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_102; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_103; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_104; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_105; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_106; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_107; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_108; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_109; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_110; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_111; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_112; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_113; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_114; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_115; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_116; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_117; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_118; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_119; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_120; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_121; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_122; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_123; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_124; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_125; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_126; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_127; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_0; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_1; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_2; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_3; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_4; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_5; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_6; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_7; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_8; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_9; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_10; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_11; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_12; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_13; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_14; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_15; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_16; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_17; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_18; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_19; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_20; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_21; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_22; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_23; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_24; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_25; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_26; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_27; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_28; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_29; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_30; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_31; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_32; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_33; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_34; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_35; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_36; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_37; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_38; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_39; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_40; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_41; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_42; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_43; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_44; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_45; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_46; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_47; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_48; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_49; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_50; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_51; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_52; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_53; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_54; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_55; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_56; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_57; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_58; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_59; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_60; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_61; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_62; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_63; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_64; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_65; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_66; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_67; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_68; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_69; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_70; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_71; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_72; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_73; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_74; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_75; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_76; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_77; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_78; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_79; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_80; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_81; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_82; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_83; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_84; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_85; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_86; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_87; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_88; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_89; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_90; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_91; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_92; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_93; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_94; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_95; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_96; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_97; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_98; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_99; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_100; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_101; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_102; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_103; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_104; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_105; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_106; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_107; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_108; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_109; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_110; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_111; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_112; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_113; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_114; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_115; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_116; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_117; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_118; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_119; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_120; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_121; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_122; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_123; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_124; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_125; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_126; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_127; // @[hh_datapath_chisel.scala 276:20]
  reg [4095:0] yj0; // @[hh_datapath_chisel.scala 53:18]
  reg [243711:0] yj_reg_1; // @[hh_datapath_chisel.scala 54:23]
  reg [243711:0] yj_reg_2; // @[hh_datapath_chisel.scala 55:23]
  reg [243711:0] yj_reg_3; // @[hh_datapath_chisel.scala 56:23]
  reg [243711:0] yj_reg_4; // @[hh_datapath_chisel.scala 57:23]
  wire [247807:0] _yj_reg_4_T_1 = {yj_reg_3[4095:0],yj_reg_4}; // @[Cat.scala 31:58]
  wire [247807:0] _yj_reg_3_T_1 = {yj_reg_2[4095:0],yj_reg_3}; // @[Cat.scala 31:58]
  wire [247807:0] _yj_reg_2_T_1 = {yj_reg_1[4095:0],yj_reg_2}; // @[Cat.scala 31:58]
  wire [247807:0] _yj_reg_1_T = {io_hh_din,yj_reg_1}; // @[Cat.scala 31:58]
  reg [4095:0] ddot_din_a_reg; // @[hh_datapath_chisel.scala 82:29]
  reg [4095:0] ddot_din_b_reg; // @[hh_datapath_chisel.scala 83:29]
  reg [4095:0] vk_reg; // @[hh_datapath_chisel.scala 85:21]
  reg [31:0] d1_reg; // @[hh_datapath_chisel.scala 86:21]
  reg [31:0] d3_reg; // @[hh_datapath_chisel.scala 87:21]
  reg [31:0] d4_update; // @[hh_datapath_chisel.scala 93:24]
  reg [31:0] x1_reg; // @[hh_datapath_chisel.scala 102:21]
  reg [31:0] d2_reg; // @[hh_datapath_chisel.scala 103:21]
  reg [31:0] vk1_reg; // @[hh_datapath_chisel.scala 104:22]
  reg [31:0] tk_reg; // @[hh_datapath_chisel.scala 105:21]
  reg [31:0] d4_reg; // @[hh_datapath_chisel.scala 106:21]
  reg [31:0] d5_reg; // @[hh_datapath_chisel.scala 107:21]
  wire [31:0] vk1_update = hqr5_io_out_s; // @[hh_datapath_chisel.scala 264:15 91:26]
  wire [31:0] vk1 = io_vk1_vld ? vk1_update : vk1_reg; // @[hh_datapath_chisel.scala 195:21 196:11 198:11]
  wire [15:0] _myNewVec_127_T_1 = io_hh_cnt + 16'h1; // @[hh_datapath_chisel.scala 234:55]
  wire [16:0] _myNewVec_127_T_2 = {{1'd0}, _myNewVec_127_T_1}; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] myVec_127 = io_hh_din[31:0]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_126 = io_hh_din[63:32]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_125 = io_hh_din[95:64]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_124 = io_hh_din[127:96]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_123 = io_hh_din[159:128]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_122 = io_hh_din[191:160]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_121 = io_hh_din[223:192]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_120 = io_hh_din[255:224]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_119 = io_hh_din[287:256]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_118 = io_hh_din[319:288]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_117 = io_hh_din[351:320]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_116 = io_hh_din[383:352]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_115 = io_hh_din[415:384]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_114 = io_hh_din[447:416]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_113 = io_hh_din[479:448]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_112 = io_hh_din[511:480]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_111 = io_hh_din[543:512]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_110 = io_hh_din[575:544]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_109 = io_hh_din[607:576]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_108 = io_hh_din[639:608]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_107 = io_hh_din[671:640]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_106 = io_hh_din[703:672]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_105 = io_hh_din[735:704]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_104 = io_hh_din[767:736]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_103 = io_hh_din[799:768]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_102 = io_hh_din[831:800]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_101 = io_hh_din[863:832]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_100 = io_hh_din[895:864]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_99 = io_hh_din[927:896]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_98 = io_hh_din[959:928]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_97 = io_hh_din[991:960]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_96 = io_hh_din[1023:992]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_95 = io_hh_din[1055:1024]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_94 = io_hh_din[1087:1056]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_93 = io_hh_din[1119:1088]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_92 = io_hh_din[1151:1120]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_91 = io_hh_din[1183:1152]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_90 = io_hh_din[1215:1184]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_89 = io_hh_din[1247:1216]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_88 = io_hh_din[1279:1248]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_87 = io_hh_din[1311:1280]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_86 = io_hh_din[1343:1312]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_85 = io_hh_din[1375:1344]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_84 = io_hh_din[1407:1376]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_83 = io_hh_din[1439:1408]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_82 = io_hh_din[1471:1440]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_81 = io_hh_din[1503:1472]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_80 = io_hh_din[1535:1504]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_79 = io_hh_din[1567:1536]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_78 = io_hh_din[1599:1568]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_77 = io_hh_din[1631:1600]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_76 = io_hh_din[1663:1632]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_75 = io_hh_din[1695:1664]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_74 = io_hh_din[1727:1696]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_73 = io_hh_din[1759:1728]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_72 = io_hh_din[1791:1760]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_71 = io_hh_din[1823:1792]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_70 = io_hh_din[1855:1824]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_69 = io_hh_din[1887:1856]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_68 = io_hh_din[1919:1888]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_67 = io_hh_din[1951:1920]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_66 = io_hh_din[1983:1952]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_65 = io_hh_din[2015:1984]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_64 = io_hh_din[2047:2016]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_63 = io_hh_din[2079:2048]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_62 = io_hh_din[2111:2080]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_61 = io_hh_din[2143:2112]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_60 = io_hh_din[2175:2144]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_59 = io_hh_din[2207:2176]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_58 = io_hh_din[2239:2208]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_57 = io_hh_din[2271:2240]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_56 = io_hh_din[2303:2272]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_55 = io_hh_din[2335:2304]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_54 = io_hh_din[2367:2336]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_53 = io_hh_din[2399:2368]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_52 = io_hh_din[2431:2400]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_51 = io_hh_din[2463:2432]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_50 = io_hh_din[2495:2464]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_49 = io_hh_din[2527:2496]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_48 = io_hh_din[2559:2528]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_47 = io_hh_din[2591:2560]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_46 = io_hh_din[2623:2592]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_45 = io_hh_din[2655:2624]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_44 = io_hh_din[2687:2656]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_43 = io_hh_din[2719:2688]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_42 = io_hh_din[2751:2720]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_41 = io_hh_din[2783:2752]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_40 = io_hh_din[2815:2784]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_39 = io_hh_din[2847:2816]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_38 = io_hh_din[2879:2848]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_37 = io_hh_din[2911:2880]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_36 = io_hh_din[2943:2912]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_35 = io_hh_din[2975:2944]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_34 = io_hh_din[3007:2976]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_33 = io_hh_din[3039:3008]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_32 = io_hh_din[3071:3040]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_31 = io_hh_din[3103:3072]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_30 = io_hh_din[3135:3104]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_29 = io_hh_din[3167:3136]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_28 = io_hh_din[3199:3168]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_27 = io_hh_din[3231:3200]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_26 = io_hh_din[3263:3232]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_25 = io_hh_din[3295:3264]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_24 = io_hh_din[3327:3296]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_23 = io_hh_din[3359:3328]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_22 = io_hh_din[3391:3360]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_21 = io_hh_din[3423:3392]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_20 = io_hh_din[3455:3424]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_19 = io_hh_din[3487:3456]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_18 = io_hh_din[3519:3488]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_17 = io_hh_din[3551:3520]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_16 = io_hh_din[3583:3552]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_15 = io_hh_din[3615:3584]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_14 = io_hh_din[3647:3616]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_13 = io_hh_din[3679:3648]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_12 = io_hh_din[3711:3680]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_11 = io_hh_din[3743:3712]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_10 = io_hh_din[3775:3744]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_9 = io_hh_din[3807:3776]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_8 = io_hh_din[3839:3808]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_7 = io_hh_din[3871:3840]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_6 = io_hh_din[3903:3872]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_5 = io_hh_din[3935:3904]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_4 = io_hh_din[3967:3936]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_3 = io_hh_din[3999:3968]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_2 = io_hh_din[4031:4000]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_1 = io_hh_din[4063:4032]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_0 = io_hh_din[4095:4064]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] _GEN_171 = 7'h1 == _myNewVec_127_T_2[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_172 = 7'h2 == _myNewVec_127_T_2[6:0] ? myVec_2 : _GEN_171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_173 = 7'h3 == _myNewVec_127_T_2[6:0] ? myVec_3 : _GEN_172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_174 = 7'h4 == _myNewVec_127_T_2[6:0] ? myVec_4 : _GEN_173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_175 = 7'h5 == _myNewVec_127_T_2[6:0] ? myVec_5 : _GEN_174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_176 = 7'h6 == _myNewVec_127_T_2[6:0] ? myVec_6 : _GEN_175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_177 = 7'h7 == _myNewVec_127_T_2[6:0] ? myVec_7 : _GEN_176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_178 = 7'h8 == _myNewVec_127_T_2[6:0] ? myVec_8 : _GEN_177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_179 = 7'h9 == _myNewVec_127_T_2[6:0] ? myVec_9 : _GEN_178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_180 = 7'ha == _myNewVec_127_T_2[6:0] ? myVec_10 : _GEN_179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_181 = 7'hb == _myNewVec_127_T_2[6:0] ? myVec_11 : _GEN_180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_182 = 7'hc == _myNewVec_127_T_2[6:0] ? myVec_12 : _GEN_181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_183 = 7'hd == _myNewVec_127_T_2[6:0] ? myVec_13 : _GEN_182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_184 = 7'he == _myNewVec_127_T_2[6:0] ? myVec_14 : _GEN_183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_185 = 7'hf == _myNewVec_127_T_2[6:0] ? myVec_15 : _GEN_184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_186 = 7'h10 == _myNewVec_127_T_2[6:0] ? myVec_16 : _GEN_185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_187 = 7'h11 == _myNewVec_127_T_2[6:0] ? myVec_17 : _GEN_186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_188 = 7'h12 == _myNewVec_127_T_2[6:0] ? myVec_18 : _GEN_187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_189 = 7'h13 == _myNewVec_127_T_2[6:0] ? myVec_19 : _GEN_188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_190 = 7'h14 == _myNewVec_127_T_2[6:0] ? myVec_20 : _GEN_189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_191 = 7'h15 == _myNewVec_127_T_2[6:0] ? myVec_21 : _GEN_190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_192 = 7'h16 == _myNewVec_127_T_2[6:0] ? myVec_22 : _GEN_191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_193 = 7'h17 == _myNewVec_127_T_2[6:0] ? myVec_23 : _GEN_192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_194 = 7'h18 == _myNewVec_127_T_2[6:0] ? myVec_24 : _GEN_193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_195 = 7'h19 == _myNewVec_127_T_2[6:0] ? myVec_25 : _GEN_194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_196 = 7'h1a == _myNewVec_127_T_2[6:0] ? myVec_26 : _GEN_195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_197 = 7'h1b == _myNewVec_127_T_2[6:0] ? myVec_27 : _GEN_196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_198 = 7'h1c == _myNewVec_127_T_2[6:0] ? myVec_28 : _GEN_197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_199 = 7'h1d == _myNewVec_127_T_2[6:0] ? myVec_29 : _GEN_198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_200 = 7'h1e == _myNewVec_127_T_2[6:0] ? myVec_30 : _GEN_199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_201 = 7'h1f == _myNewVec_127_T_2[6:0] ? myVec_31 : _GEN_200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_202 = 7'h20 == _myNewVec_127_T_2[6:0] ? myVec_32 : _GEN_201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_203 = 7'h21 == _myNewVec_127_T_2[6:0] ? myVec_33 : _GEN_202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_204 = 7'h22 == _myNewVec_127_T_2[6:0] ? myVec_34 : _GEN_203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_205 = 7'h23 == _myNewVec_127_T_2[6:0] ? myVec_35 : _GEN_204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_206 = 7'h24 == _myNewVec_127_T_2[6:0] ? myVec_36 : _GEN_205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_207 = 7'h25 == _myNewVec_127_T_2[6:0] ? myVec_37 : _GEN_206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_208 = 7'h26 == _myNewVec_127_T_2[6:0] ? myVec_38 : _GEN_207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_209 = 7'h27 == _myNewVec_127_T_2[6:0] ? myVec_39 : _GEN_208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_210 = 7'h28 == _myNewVec_127_T_2[6:0] ? myVec_40 : _GEN_209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_211 = 7'h29 == _myNewVec_127_T_2[6:0] ? myVec_41 : _GEN_210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_212 = 7'h2a == _myNewVec_127_T_2[6:0] ? myVec_42 : _GEN_211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_213 = 7'h2b == _myNewVec_127_T_2[6:0] ? myVec_43 : _GEN_212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_214 = 7'h2c == _myNewVec_127_T_2[6:0] ? myVec_44 : _GEN_213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_215 = 7'h2d == _myNewVec_127_T_2[6:0] ? myVec_45 : _GEN_214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_216 = 7'h2e == _myNewVec_127_T_2[6:0] ? myVec_46 : _GEN_215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_217 = 7'h2f == _myNewVec_127_T_2[6:0] ? myVec_47 : _GEN_216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_218 = 7'h30 == _myNewVec_127_T_2[6:0] ? myVec_48 : _GEN_217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_219 = 7'h31 == _myNewVec_127_T_2[6:0] ? myVec_49 : _GEN_218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_220 = 7'h32 == _myNewVec_127_T_2[6:0] ? myVec_50 : _GEN_219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_221 = 7'h33 == _myNewVec_127_T_2[6:0] ? myVec_51 : _GEN_220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_222 = 7'h34 == _myNewVec_127_T_2[6:0] ? myVec_52 : _GEN_221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_223 = 7'h35 == _myNewVec_127_T_2[6:0] ? myVec_53 : _GEN_222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_224 = 7'h36 == _myNewVec_127_T_2[6:0] ? myVec_54 : _GEN_223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_225 = 7'h37 == _myNewVec_127_T_2[6:0] ? myVec_55 : _GEN_224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_226 = 7'h38 == _myNewVec_127_T_2[6:0] ? myVec_56 : _GEN_225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_227 = 7'h39 == _myNewVec_127_T_2[6:0] ? myVec_57 : _GEN_226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_228 = 7'h3a == _myNewVec_127_T_2[6:0] ? myVec_58 : _GEN_227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_229 = 7'h3b == _myNewVec_127_T_2[6:0] ? myVec_59 : _GEN_228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_230 = 7'h3c == _myNewVec_127_T_2[6:0] ? myVec_60 : _GEN_229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_231 = 7'h3d == _myNewVec_127_T_2[6:0] ? myVec_61 : _GEN_230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_232 = 7'h3e == _myNewVec_127_T_2[6:0] ? myVec_62 : _GEN_231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_233 = 7'h3f == _myNewVec_127_T_2[6:0] ? myVec_63 : _GEN_232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_234 = 7'h40 == _myNewVec_127_T_2[6:0] ? myVec_64 : _GEN_233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_235 = 7'h41 == _myNewVec_127_T_2[6:0] ? myVec_65 : _GEN_234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_236 = 7'h42 == _myNewVec_127_T_2[6:0] ? myVec_66 : _GEN_235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_237 = 7'h43 == _myNewVec_127_T_2[6:0] ? myVec_67 : _GEN_236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_238 = 7'h44 == _myNewVec_127_T_2[6:0] ? myVec_68 : _GEN_237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_239 = 7'h45 == _myNewVec_127_T_2[6:0] ? myVec_69 : _GEN_238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_240 = 7'h46 == _myNewVec_127_T_2[6:0] ? myVec_70 : _GEN_239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_241 = 7'h47 == _myNewVec_127_T_2[6:0] ? myVec_71 : _GEN_240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_242 = 7'h48 == _myNewVec_127_T_2[6:0] ? myVec_72 : _GEN_241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_243 = 7'h49 == _myNewVec_127_T_2[6:0] ? myVec_73 : _GEN_242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_244 = 7'h4a == _myNewVec_127_T_2[6:0] ? myVec_74 : _GEN_243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_245 = 7'h4b == _myNewVec_127_T_2[6:0] ? myVec_75 : _GEN_244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_246 = 7'h4c == _myNewVec_127_T_2[6:0] ? myVec_76 : _GEN_245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_247 = 7'h4d == _myNewVec_127_T_2[6:0] ? myVec_77 : _GEN_246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_248 = 7'h4e == _myNewVec_127_T_2[6:0] ? myVec_78 : _GEN_247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_249 = 7'h4f == _myNewVec_127_T_2[6:0] ? myVec_79 : _GEN_248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_250 = 7'h50 == _myNewVec_127_T_2[6:0] ? myVec_80 : _GEN_249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_251 = 7'h51 == _myNewVec_127_T_2[6:0] ? myVec_81 : _GEN_250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_252 = 7'h52 == _myNewVec_127_T_2[6:0] ? myVec_82 : _GEN_251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_253 = 7'h53 == _myNewVec_127_T_2[6:0] ? myVec_83 : _GEN_252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_254 = 7'h54 == _myNewVec_127_T_2[6:0] ? myVec_84 : _GEN_253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_255 = 7'h55 == _myNewVec_127_T_2[6:0] ? myVec_85 : _GEN_254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_256 = 7'h56 == _myNewVec_127_T_2[6:0] ? myVec_86 : _GEN_255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_257 = 7'h57 == _myNewVec_127_T_2[6:0] ? myVec_87 : _GEN_256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_258 = 7'h58 == _myNewVec_127_T_2[6:0] ? myVec_88 : _GEN_257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_259 = 7'h59 == _myNewVec_127_T_2[6:0] ? myVec_89 : _GEN_258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_260 = 7'h5a == _myNewVec_127_T_2[6:0] ? myVec_90 : _GEN_259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_261 = 7'h5b == _myNewVec_127_T_2[6:0] ? myVec_91 : _GEN_260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_262 = 7'h5c == _myNewVec_127_T_2[6:0] ? myVec_92 : _GEN_261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_263 = 7'h5d == _myNewVec_127_T_2[6:0] ? myVec_93 : _GEN_262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_264 = 7'h5e == _myNewVec_127_T_2[6:0] ? myVec_94 : _GEN_263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_265 = 7'h5f == _myNewVec_127_T_2[6:0] ? myVec_95 : _GEN_264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_266 = 7'h60 == _myNewVec_127_T_2[6:0] ? myVec_96 : _GEN_265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_267 = 7'h61 == _myNewVec_127_T_2[6:0] ? myVec_97 : _GEN_266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_268 = 7'h62 == _myNewVec_127_T_2[6:0] ? myVec_98 : _GEN_267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_269 = 7'h63 == _myNewVec_127_T_2[6:0] ? myVec_99 : _GEN_268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_270 = 7'h64 == _myNewVec_127_T_2[6:0] ? myVec_100 : _GEN_269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_271 = 7'h65 == _myNewVec_127_T_2[6:0] ? myVec_101 : _GEN_270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_272 = 7'h66 == _myNewVec_127_T_2[6:0] ? myVec_102 : _GEN_271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_273 = 7'h67 == _myNewVec_127_T_2[6:0] ? myVec_103 : _GEN_272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_274 = 7'h68 == _myNewVec_127_T_2[6:0] ? myVec_104 : _GEN_273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_275 = 7'h69 == _myNewVec_127_T_2[6:0] ? myVec_105 : _GEN_274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_276 = 7'h6a == _myNewVec_127_T_2[6:0] ? myVec_106 : _GEN_275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_277 = 7'h6b == _myNewVec_127_T_2[6:0] ? myVec_107 : _GEN_276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_278 = 7'h6c == _myNewVec_127_T_2[6:0] ? myVec_108 : _GEN_277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_279 = 7'h6d == _myNewVec_127_T_2[6:0] ? myVec_109 : _GEN_278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_280 = 7'h6e == _myNewVec_127_T_2[6:0] ? myVec_110 : _GEN_279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_281 = 7'h6f == _myNewVec_127_T_2[6:0] ? myVec_111 : _GEN_280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_282 = 7'h70 == _myNewVec_127_T_2[6:0] ? myVec_112 : _GEN_281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_283 = 7'h71 == _myNewVec_127_T_2[6:0] ? myVec_113 : _GEN_282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_284 = 7'h72 == _myNewVec_127_T_2[6:0] ? myVec_114 : _GEN_283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_285 = 7'h73 == _myNewVec_127_T_2[6:0] ? myVec_115 : _GEN_284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_286 = 7'h74 == _myNewVec_127_T_2[6:0] ? myVec_116 : _GEN_285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_287 = 7'h75 == _myNewVec_127_T_2[6:0] ? myVec_117 : _GEN_286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_288 = 7'h76 == _myNewVec_127_T_2[6:0] ? myVec_118 : _GEN_287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_289 = 7'h77 == _myNewVec_127_T_2[6:0] ? myVec_119 : _GEN_288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_290 = 7'h78 == _myNewVec_127_T_2[6:0] ? myVec_120 : _GEN_289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_291 = 7'h79 == _myNewVec_127_T_2[6:0] ? myVec_121 : _GEN_290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_292 = 7'h7a == _myNewVec_127_T_2[6:0] ? myVec_122 : _GEN_291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_293 = 7'h7b == _myNewVec_127_T_2[6:0] ? myVec_123 : _GEN_292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_294 = 7'h7c == _myNewVec_127_T_2[6:0] ? myVec_124 : _GEN_293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_295 = 7'h7d == _myNewVec_127_T_2[6:0] ? myVec_125 : _GEN_294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_296 = 7'h7e == _myNewVec_127_T_2[6:0] ? myVec_126 : _GEN_295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_127 = 7'h7f == _myNewVec_127_T_2[6:0] ? myVec_127 : _GEN_296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_126_T_3 = _myNewVec_127_T_1 + 16'h1; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_299 = 7'h1 == _myNewVec_126_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_300 = 7'h2 == _myNewVec_126_T_3[6:0] ? myVec_2 : _GEN_299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_301 = 7'h3 == _myNewVec_126_T_3[6:0] ? myVec_3 : _GEN_300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_302 = 7'h4 == _myNewVec_126_T_3[6:0] ? myVec_4 : _GEN_301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_303 = 7'h5 == _myNewVec_126_T_3[6:0] ? myVec_5 : _GEN_302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_304 = 7'h6 == _myNewVec_126_T_3[6:0] ? myVec_6 : _GEN_303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_305 = 7'h7 == _myNewVec_126_T_3[6:0] ? myVec_7 : _GEN_304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_306 = 7'h8 == _myNewVec_126_T_3[6:0] ? myVec_8 : _GEN_305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_307 = 7'h9 == _myNewVec_126_T_3[6:0] ? myVec_9 : _GEN_306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_308 = 7'ha == _myNewVec_126_T_3[6:0] ? myVec_10 : _GEN_307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_309 = 7'hb == _myNewVec_126_T_3[6:0] ? myVec_11 : _GEN_308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_310 = 7'hc == _myNewVec_126_T_3[6:0] ? myVec_12 : _GEN_309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_311 = 7'hd == _myNewVec_126_T_3[6:0] ? myVec_13 : _GEN_310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_312 = 7'he == _myNewVec_126_T_3[6:0] ? myVec_14 : _GEN_311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_313 = 7'hf == _myNewVec_126_T_3[6:0] ? myVec_15 : _GEN_312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_314 = 7'h10 == _myNewVec_126_T_3[6:0] ? myVec_16 : _GEN_313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_315 = 7'h11 == _myNewVec_126_T_3[6:0] ? myVec_17 : _GEN_314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_316 = 7'h12 == _myNewVec_126_T_3[6:0] ? myVec_18 : _GEN_315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_317 = 7'h13 == _myNewVec_126_T_3[6:0] ? myVec_19 : _GEN_316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_318 = 7'h14 == _myNewVec_126_T_3[6:0] ? myVec_20 : _GEN_317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_319 = 7'h15 == _myNewVec_126_T_3[6:0] ? myVec_21 : _GEN_318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_320 = 7'h16 == _myNewVec_126_T_3[6:0] ? myVec_22 : _GEN_319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_321 = 7'h17 == _myNewVec_126_T_3[6:0] ? myVec_23 : _GEN_320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_322 = 7'h18 == _myNewVec_126_T_3[6:0] ? myVec_24 : _GEN_321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_323 = 7'h19 == _myNewVec_126_T_3[6:0] ? myVec_25 : _GEN_322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_324 = 7'h1a == _myNewVec_126_T_3[6:0] ? myVec_26 : _GEN_323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_325 = 7'h1b == _myNewVec_126_T_3[6:0] ? myVec_27 : _GEN_324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_326 = 7'h1c == _myNewVec_126_T_3[6:0] ? myVec_28 : _GEN_325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_327 = 7'h1d == _myNewVec_126_T_3[6:0] ? myVec_29 : _GEN_326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_328 = 7'h1e == _myNewVec_126_T_3[6:0] ? myVec_30 : _GEN_327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_329 = 7'h1f == _myNewVec_126_T_3[6:0] ? myVec_31 : _GEN_328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_330 = 7'h20 == _myNewVec_126_T_3[6:0] ? myVec_32 : _GEN_329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_331 = 7'h21 == _myNewVec_126_T_3[6:0] ? myVec_33 : _GEN_330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_332 = 7'h22 == _myNewVec_126_T_3[6:0] ? myVec_34 : _GEN_331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_333 = 7'h23 == _myNewVec_126_T_3[6:0] ? myVec_35 : _GEN_332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_334 = 7'h24 == _myNewVec_126_T_3[6:0] ? myVec_36 : _GEN_333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_335 = 7'h25 == _myNewVec_126_T_3[6:0] ? myVec_37 : _GEN_334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_336 = 7'h26 == _myNewVec_126_T_3[6:0] ? myVec_38 : _GEN_335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_337 = 7'h27 == _myNewVec_126_T_3[6:0] ? myVec_39 : _GEN_336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_338 = 7'h28 == _myNewVec_126_T_3[6:0] ? myVec_40 : _GEN_337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_339 = 7'h29 == _myNewVec_126_T_3[6:0] ? myVec_41 : _GEN_338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_340 = 7'h2a == _myNewVec_126_T_3[6:0] ? myVec_42 : _GEN_339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_341 = 7'h2b == _myNewVec_126_T_3[6:0] ? myVec_43 : _GEN_340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_342 = 7'h2c == _myNewVec_126_T_3[6:0] ? myVec_44 : _GEN_341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_343 = 7'h2d == _myNewVec_126_T_3[6:0] ? myVec_45 : _GEN_342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_344 = 7'h2e == _myNewVec_126_T_3[6:0] ? myVec_46 : _GEN_343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_345 = 7'h2f == _myNewVec_126_T_3[6:0] ? myVec_47 : _GEN_344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_346 = 7'h30 == _myNewVec_126_T_3[6:0] ? myVec_48 : _GEN_345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_347 = 7'h31 == _myNewVec_126_T_3[6:0] ? myVec_49 : _GEN_346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_348 = 7'h32 == _myNewVec_126_T_3[6:0] ? myVec_50 : _GEN_347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_349 = 7'h33 == _myNewVec_126_T_3[6:0] ? myVec_51 : _GEN_348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_350 = 7'h34 == _myNewVec_126_T_3[6:0] ? myVec_52 : _GEN_349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_351 = 7'h35 == _myNewVec_126_T_3[6:0] ? myVec_53 : _GEN_350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_352 = 7'h36 == _myNewVec_126_T_3[6:0] ? myVec_54 : _GEN_351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_353 = 7'h37 == _myNewVec_126_T_3[6:0] ? myVec_55 : _GEN_352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_354 = 7'h38 == _myNewVec_126_T_3[6:0] ? myVec_56 : _GEN_353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_355 = 7'h39 == _myNewVec_126_T_3[6:0] ? myVec_57 : _GEN_354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_356 = 7'h3a == _myNewVec_126_T_3[6:0] ? myVec_58 : _GEN_355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_357 = 7'h3b == _myNewVec_126_T_3[6:0] ? myVec_59 : _GEN_356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_358 = 7'h3c == _myNewVec_126_T_3[6:0] ? myVec_60 : _GEN_357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_359 = 7'h3d == _myNewVec_126_T_3[6:0] ? myVec_61 : _GEN_358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_360 = 7'h3e == _myNewVec_126_T_3[6:0] ? myVec_62 : _GEN_359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_361 = 7'h3f == _myNewVec_126_T_3[6:0] ? myVec_63 : _GEN_360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_362 = 7'h40 == _myNewVec_126_T_3[6:0] ? myVec_64 : _GEN_361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_363 = 7'h41 == _myNewVec_126_T_3[6:0] ? myVec_65 : _GEN_362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_364 = 7'h42 == _myNewVec_126_T_3[6:0] ? myVec_66 : _GEN_363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_365 = 7'h43 == _myNewVec_126_T_3[6:0] ? myVec_67 : _GEN_364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_366 = 7'h44 == _myNewVec_126_T_3[6:0] ? myVec_68 : _GEN_365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_367 = 7'h45 == _myNewVec_126_T_3[6:0] ? myVec_69 : _GEN_366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_368 = 7'h46 == _myNewVec_126_T_3[6:0] ? myVec_70 : _GEN_367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_369 = 7'h47 == _myNewVec_126_T_3[6:0] ? myVec_71 : _GEN_368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_370 = 7'h48 == _myNewVec_126_T_3[6:0] ? myVec_72 : _GEN_369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_371 = 7'h49 == _myNewVec_126_T_3[6:0] ? myVec_73 : _GEN_370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_372 = 7'h4a == _myNewVec_126_T_3[6:0] ? myVec_74 : _GEN_371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_373 = 7'h4b == _myNewVec_126_T_3[6:0] ? myVec_75 : _GEN_372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_374 = 7'h4c == _myNewVec_126_T_3[6:0] ? myVec_76 : _GEN_373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_375 = 7'h4d == _myNewVec_126_T_3[6:0] ? myVec_77 : _GEN_374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_376 = 7'h4e == _myNewVec_126_T_3[6:0] ? myVec_78 : _GEN_375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_377 = 7'h4f == _myNewVec_126_T_3[6:0] ? myVec_79 : _GEN_376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_378 = 7'h50 == _myNewVec_126_T_3[6:0] ? myVec_80 : _GEN_377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_379 = 7'h51 == _myNewVec_126_T_3[6:0] ? myVec_81 : _GEN_378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_380 = 7'h52 == _myNewVec_126_T_3[6:0] ? myVec_82 : _GEN_379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_381 = 7'h53 == _myNewVec_126_T_3[6:0] ? myVec_83 : _GEN_380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_382 = 7'h54 == _myNewVec_126_T_3[6:0] ? myVec_84 : _GEN_381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_383 = 7'h55 == _myNewVec_126_T_3[6:0] ? myVec_85 : _GEN_382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_384 = 7'h56 == _myNewVec_126_T_3[6:0] ? myVec_86 : _GEN_383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_385 = 7'h57 == _myNewVec_126_T_3[6:0] ? myVec_87 : _GEN_384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_386 = 7'h58 == _myNewVec_126_T_3[6:0] ? myVec_88 : _GEN_385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_387 = 7'h59 == _myNewVec_126_T_3[6:0] ? myVec_89 : _GEN_386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_388 = 7'h5a == _myNewVec_126_T_3[6:0] ? myVec_90 : _GEN_387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_389 = 7'h5b == _myNewVec_126_T_3[6:0] ? myVec_91 : _GEN_388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_390 = 7'h5c == _myNewVec_126_T_3[6:0] ? myVec_92 : _GEN_389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_391 = 7'h5d == _myNewVec_126_T_3[6:0] ? myVec_93 : _GEN_390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_392 = 7'h5e == _myNewVec_126_T_3[6:0] ? myVec_94 : _GEN_391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_393 = 7'h5f == _myNewVec_126_T_3[6:0] ? myVec_95 : _GEN_392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_394 = 7'h60 == _myNewVec_126_T_3[6:0] ? myVec_96 : _GEN_393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_395 = 7'h61 == _myNewVec_126_T_3[6:0] ? myVec_97 : _GEN_394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_396 = 7'h62 == _myNewVec_126_T_3[6:0] ? myVec_98 : _GEN_395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_397 = 7'h63 == _myNewVec_126_T_3[6:0] ? myVec_99 : _GEN_396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_398 = 7'h64 == _myNewVec_126_T_3[6:0] ? myVec_100 : _GEN_397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_399 = 7'h65 == _myNewVec_126_T_3[6:0] ? myVec_101 : _GEN_398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_400 = 7'h66 == _myNewVec_126_T_3[6:0] ? myVec_102 : _GEN_399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_401 = 7'h67 == _myNewVec_126_T_3[6:0] ? myVec_103 : _GEN_400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_402 = 7'h68 == _myNewVec_126_T_3[6:0] ? myVec_104 : _GEN_401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_403 = 7'h69 == _myNewVec_126_T_3[6:0] ? myVec_105 : _GEN_402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_404 = 7'h6a == _myNewVec_126_T_3[6:0] ? myVec_106 : _GEN_403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_405 = 7'h6b == _myNewVec_126_T_3[6:0] ? myVec_107 : _GEN_404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_406 = 7'h6c == _myNewVec_126_T_3[6:0] ? myVec_108 : _GEN_405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_407 = 7'h6d == _myNewVec_126_T_3[6:0] ? myVec_109 : _GEN_406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_408 = 7'h6e == _myNewVec_126_T_3[6:0] ? myVec_110 : _GEN_407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_409 = 7'h6f == _myNewVec_126_T_3[6:0] ? myVec_111 : _GEN_408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_410 = 7'h70 == _myNewVec_126_T_3[6:0] ? myVec_112 : _GEN_409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_411 = 7'h71 == _myNewVec_126_T_3[6:0] ? myVec_113 : _GEN_410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_412 = 7'h72 == _myNewVec_126_T_3[6:0] ? myVec_114 : _GEN_411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_413 = 7'h73 == _myNewVec_126_T_3[6:0] ? myVec_115 : _GEN_412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_414 = 7'h74 == _myNewVec_126_T_3[6:0] ? myVec_116 : _GEN_413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_415 = 7'h75 == _myNewVec_126_T_3[6:0] ? myVec_117 : _GEN_414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_416 = 7'h76 == _myNewVec_126_T_3[6:0] ? myVec_118 : _GEN_415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_417 = 7'h77 == _myNewVec_126_T_3[6:0] ? myVec_119 : _GEN_416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_418 = 7'h78 == _myNewVec_126_T_3[6:0] ? myVec_120 : _GEN_417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_419 = 7'h79 == _myNewVec_126_T_3[6:0] ? myVec_121 : _GEN_418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_420 = 7'h7a == _myNewVec_126_T_3[6:0] ? myVec_122 : _GEN_419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_421 = 7'h7b == _myNewVec_126_T_3[6:0] ? myVec_123 : _GEN_420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_422 = 7'h7c == _myNewVec_126_T_3[6:0] ? myVec_124 : _GEN_421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_423 = 7'h7d == _myNewVec_126_T_3[6:0] ? myVec_125 : _GEN_422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_424 = 7'h7e == _myNewVec_126_T_3[6:0] ? myVec_126 : _GEN_423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_126 = 7'h7f == _myNewVec_126_T_3[6:0] ? myVec_127 : _GEN_424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_125_T_3 = _myNewVec_127_T_1 + 16'h2; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_427 = 7'h1 == _myNewVec_125_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_428 = 7'h2 == _myNewVec_125_T_3[6:0] ? myVec_2 : _GEN_427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_429 = 7'h3 == _myNewVec_125_T_3[6:0] ? myVec_3 : _GEN_428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_430 = 7'h4 == _myNewVec_125_T_3[6:0] ? myVec_4 : _GEN_429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_431 = 7'h5 == _myNewVec_125_T_3[6:0] ? myVec_5 : _GEN_430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_432 = 7'h6 == _myNewVec_125_T_3[6:0] ? myVec_6 : _GEN_431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_433 = 7'h7 == _myNewVec_125_T_3[6:0] ? myVec_7 : _GEN_432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_434 = 7'h8 == _myNewVec_125_T_3[6:0] ? myVec_8 : _GEN_433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_435 = 7'h9 == _myNewVec_125_T_3[6:0] ? myVec_9 : _GEN_434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_436 = 7'ha == _myNewVec_125_T_3[6:0] ? myVec_10 : _GEN_435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_437 = 7'hb == _myNewVec_125_T_3[6:0] ? myVec_11 : _GEN_436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_438 = 7'hc == _myNewVec_125_T_3[6:0] ? myVec_12 : _GEN_437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_439 = 7'hd == _myNewVec_125_T_3[6:0] ? myVec_13 : _GEN_438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_440 = 7'he == _myNewVec_125_T_3[6:0] ? myVec_14 : _GEN_439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_441 = 7'hf == _myNewVec_125_T_3[6:0] ? myVec_15 : _GEN_440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_442 = 7'h10 == _myNewVec_125_T_3[6:0] ? myVec_16 : _GEN_441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_443 = 7'h11 == _myNewVec_125_T_3[6:0] ? myVec_17 : _GEN_442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_444 = 7'h12 == _myNewVec_125_T_3[6:0] ? myVec_18 : _GEN_443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_445 = 7'h13 == _myNewVec_125_T_3[6:0] ? myVec_19 : _GEN_444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_446 = 7'h14 == _myNewVec_125_T_3[6:0] ? myVec_20 : _GEN_445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_447 = 7'h15 == _myNewVec_125_T_3[6:0] ? myVec_21 : _GEN_446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_448 = 7'h16 == _myNewVec_125_T_3[6:0] ? myVec_22 : _GEN_447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_449 = 7'h17 == _myNewVec_125_T_3[6:0] ? myVec_23 : _GEN_448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_450 = 7'h18 == _myNewVec_125_T_3[6:0] ? myVec_24 : _GEN_449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_451 = 7'h19 == _myNewVec_125_T_3[6:0] ? myVec_25 : _GEN_450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_452 = 7'h1a == _myNewVec_125_T_3[6:0] ? myVec_26 : _GEN_451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_453 = 7'h1b == _myNewVec_125_T_3[6:0] ? myVec_27 : _GEN_452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_454 = 7'h1c == _myNewVec_125_T_3[6:0] ? myVec_28 : _GEN_453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_455 = 7'h1d == _myNewVec_125_T_3[6:0] ? myVec_29 : _GEN_454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_456 = 7'h1e == _myNewVec_125_T_3[6:0] ? myVec_30 : _GEN_455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_457 = 7'h1f == _myNewVec_125_T_3[6:0] ? myVec_31 : _GEN_456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_458 = 7'h20 == _myNewVec_125_T_3[6:0] ? myVec_32 : _GEN_457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_459 = 7'h21 == _myNewVec_125_T_3[6:0] ? myVec_33 : _GEN_458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_460 = 7'h22 == _myNewVec_125_T_3[6:0] ? myVec_34 : _GEN_459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_461 = 7'h23 == _myNewVec_125_T_3[6:0] ? myVec_35 : _GEN_460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_462 = 7'h24 == _myNewVec_125_T_3[6:0] ? myVec_36 : _GEN_461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_463 = 7'h25 == _myNewVec_125_T_3[6:0] ? myVec_37 : _GEN_462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_464 = 7'h26 == _myNewVec_125_T_3[6:0] ? myVec_38 : _GEN_463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_465 = 7'h27 == _myNewVec_125_T_3[6:0] ? myVec_39 : _GEN_464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_466 = 7'h28 == _myNewVec_125_T_3[6:0] ? myVec_40 : _GEN_465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_467 = 7'h29 == _myNewVec_125_T_3[6:0] ? myVec_41 : _GEN_466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_468 = 7'h2a == _myNewVec_125_T_3[6:0] ? myVec_42 : _GEN_467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_469 = 7'h2b == _myNewVec_125_T_3[6:0] ? myVec_43 : _GEN_468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_470 = 7'h2c == _myNewVec_125_T_3[6:0] ? myVec_44 : _GEN_469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_471 = 7'h2d == _myNewVec_125_T_3[6:0] ? myVec_45 : _GEN_470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_472 = 7'h2e == _myNewVec_125_T_3[6:0] ? myVec_46 : _GEN_471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_473 = 7'h2f == _myNewVec_125_T_3[6:0] ? myVec_47 : _GEN_472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_474 = 7'h30 == _myNewVec_125_T_3[6:0] ? myVec_48 : _GEN_473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_475 = 7'h31 == _myNewVec_125_T_3[6:0] ? myVec_49 : _GEN_474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_476 = 7'h32 == _myNewVec_125_T_3[6:0] ? myVec_50 : _GEN_475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_477 = 7'h33 == _myNewVec_125_T_3[6:0] ? myVec_51 : _GEN_476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_478 = 7'h34 == _myNewVec_125_T_3[6:0] ? myVec_52 : _GEN_477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_479 = 7'h35 == _myNewVec_125_T_3[6:0] ? myVec_53 : _GEN_478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_480 = 7'h36 == _myNewVec_125_T_3[6:0] ? myVec_54 : _GEN_479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_481 = 7'h37 == _myNewVec_125_T_3[6:0] ? myVec_55 : _GEN_480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_482 = 7'h38 == _myNewVec_125_T_3[6:0] ? myVec_56 : _GEN_481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_483 = 7'h39 == _myNewVec_125_T_3[6:0] ? myVec_57 : _GEN_482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_484 = 7'h3a == _myNewVec_125_T_3[6:0] ? myVec_58 : _GEN_483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_485 = 7'h3b == _myNewVec_125_T_3[6:0] ? myVec_59 : _GEN_484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_486 = 7'h3c == _myNewVec_125_T_3[6:0] ? myVec_60 : _GEN_485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_487 = 7'h3d == _myNewVec_125_T_3[6:0] ? myVec_61 : _GEN_486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_488 = 7'h3e == _myNewVec_125_T_3[6:0] ? myVec_62 : _GEN_487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_489 = 7'h3f == _myNewVec_125_T_3[6:0] ? myVec_63 : _GEN_488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_490 = 7'h40 == _myNewVec_125_T_3[6:0] ? myVec_64 : _GEN_489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_491 = 7'h41 == _myNewVec_125_T_3[6:0] ? myVec_65 : _GEN_490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_492 = 7'h42 == _myNewVec_125_T_3[6:0] ? myVec_66 : _GEN_491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_493 = 7'h43 == _myNewVec_125_T_3[6:0] ? myVec_67 : _GEN_492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_494 = 7'h44 == _myNewVec_125_T_3[6:0] ? myVec_68 : _GEN_493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_495 = 7'h45 == _myNewVec_125_T_3[6:0] ? myVec_69 : _GEN_494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_496 = 7'h46 == _myNewVec_125_T_3[6:0] ? myVec_70 : _GEN_495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_497 = 7'h47 == _myNewVec_125_T_3[6:0] ? myVec_71 : _GEN_496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_498 = 7'h48 == _myNewVec_125_T_3[6:0] ? myVec_72 : _GEN_497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_499 = 7'h49 == _myNewVec_125_T_3[6:0] ? myVec_73 : _GEN_498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_500 = 7'h4a == _myNewVec_125_T_3[6:0] ? myVec_74 : _GEN_499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_501 = 7'h4b == _myNewVec_125_T_3[6:0] ? myVec_75 : _GEN_500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_502 = 7'h4c == _myNewVec_125_T_3[6:0] ? myVec_76 : _GEN_501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_503 = 7'h4d == _myNewVec_125_T_3[6:0] ? myVec_77 : _GEN_502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_504 = 7'h4e == _myNewVec_125_T_3[6:0] ? myVec_78 : _GEN_503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_505 = 7'h4f == _myNewVec_125_T_3[6:0] ? myVec_79 : _GEN_504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_506 = 7'h50 == _myNewVec_125_T_3[6:0] ? myVec_80 : _GEN_505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_507 = 7'h51 == _myNewVec_125_T_3[6:0] ? myVec_81 : _GEN_506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_508 = 7'h52 == _myNewVec_125_T_3[6:0] ? myVec_82 : _GEN_507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_509 = 7'h53 == _myNewVec_125_T_3[6:0] ? myVec_83 : _GEN_508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_510 = 7'h54 == _myNewVec_125_T_3[6:0] ? myVec_84 : _GEN_509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_511 = 7'h55 == _myNewVec_125_T_3[6:0] ? myVec_85 : _GEN_510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_512 = 7'h56 == _myNewVec_125_T_3[6:0] ? myVec_86 : _GEN_511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_513 = 7'h57 == _myNewVec_125_T_3[6:0] ? myVec_87 : _GEN_512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_514 = 7'h58 == _myNewVec_125_T_3[6:0] ? myVec_88 : _GEN_513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_515 = 7'h59 == _myNewVec_125_T_3[6:0] ? myVec_89 : _GEN_514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_516 = 7'h5a == _myNewVec_125_T_3[6:0] ? myVec_90 : _GEN_515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_517 = 7'h5b == _myNewVec_125_T_3[6:0] ? myVec_91 : _GEN_516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_518 = 7'h5c == _myNewVec_125_T_3[6:0] ? myVec_92 : _GEN_517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_519 = 7'h5d == _myNewVec_125_T_3[6:0] ? myVec_93 : _GEN_518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_520 = 7'h5e == _myNewVec_125_T_3[6:0] ? myVec_94 : _GEN_519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_521 = 7'h5f == _myNewVec_125_T_3[6:0] ? myVec_95 : _GEN_520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_522 = 7'h60 == _myNewVec_125_T_3[6:0] ? myVec_96 : _GEN_521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_523 = 7'h61 == _myNewVec_125_T_3[6:0] ? myVec_97 : _GEN_522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_524 = 7'h62 == _myNewVec_125_T_3[6:0] ? myVec_98 : _GEN_523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_525 = 7'h63 == _myNewVec_125_T_3[6:0] ? myVec_99 : _GEN_524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_526 = 7'h64 == _myNewVec_125_T_3[6:0] ? myVec_100 : _GEN_525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_527 = 7'h65 == _myNewVec_125_T_3[6:0] ? myVec_101 : _GEN_526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_528 = 7'h66 == _myNewVec_125_T_3[6:0] ? myVec_102 : _GEN_527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_529 = 7'h67 == _myNewVec_125_T_3[6:0] ? myVec_103 : _GEN_528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_530 = 7'h68 == _myNewVec_125_T_3[6:0] ? myVec_104 : _GEN_529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_531 = 7'h69 == _myNewVec_125_T_3[6:0] ? myVec_105 : _GEN_530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_532 = 7'h6a == _myNewVec_125_T_3[6:0] ? myVec_106 : _GEN_531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_533 = 7'h6b == _myNewVec_125_T_3[6:0] ? myVec_107 : _GEN_532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_534 = 7'h6c == _myNewVec_125_T_3[6:0] ? myVec_108 : _GEN_533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_535 = 7'h6d == _myNewVec_125_T_3[6:0] ? myVec_109 : _GEN_534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_536 = 7'h6e == _myNewVec_125_T_3[6:0] ? myVec_110 : _GEN_535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_537 = 7'h6f == _myNewVec_125_T_3[6:0] ? myVec_111 : _GEN_536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_538 = 7'h70 == _myNewVec_125_T_3[6:0] ? myVec_112 : _GEN_537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_539 = 7'h71 == _myNewVec_125_T_3[6:0] ? myVec_113 : _GEN_538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_540 = 7'h72 == _myNewVec_125_T_3[6:0] ? myVec_114 : _GEN_539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_541 = 7'h73 == _myNewVec_125_T_3[6:0] ? myVec_115 : _GEN_540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_542 = 7'h74 == _myNewVec_125_T_3[6:0] ? myVec_116 : _GEN_541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_543 = 7'h75 == _myNewVec_125_T_3[6:0] ? myVec_117 : _GEN_542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_544 = 7'h76 == _myNewVec_125_T_3[6:0] ? myVec_118 : _GEN_543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_545 = 7'h77 == _myNewVec_125_T_3[6:0] ? myVec_119 : _GEN_544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_546 = 7'h78 == _myNewVec_125_T_3[6:0] ? myVec_120 : _GEN_545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_547 = 7'h79 == _myNewVec_125_T_3[6:0] ? myVec_121 : _GEN_546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_548 = 7'h7a == _myNewVec_125_T_3[6:0] ? myVec_122 : _GEN_547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_549 = 7'h7b == _myNewVec_125_T_3[6:0] ? myVec_123 : _GEN_548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_550 = 7'h7c == _myNewVec_125_T_3[6:0] ? myVec_124 : _GEN_549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_551 = 7'h7d == _myNewVec_125_T_3[6:0] ? myVec_125 : _GEN_550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_552 = 7'h7e == _myNewVec_125_T_3[6:0] ? myVec_126 : _GEN_551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_125 = 7'h7f == _myNewVec_125_T_3[6:0] ? myVec_127 : _GEN_552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_124_T_3 = _myNewVec_127_T_1 + 16'h3; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_555 = 7'h1 == _myNewVec_124_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_556 = 7'h2 == _myNewVec_124_T_3[6:0] ? myVec_2 : _GEN_555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_557 = 7'h3 == _myNewVec_124_T_3[6:0] ? myVec_3 : _GEN_556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_558 = 7'h4 == _myNewVec_124_T_3[6:0] ? myVec_4 : _GEN_557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_559 = 7'h5 == _myNewVec_124_T_3[6:0] ? myVec_5 : _GEN_558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_560 = 7'h6 == _myNewVec_124_T_3[6:0] ? myVec_6 : _GEN_559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_561 = 7'h7 == _myNewVec_124_T_3[6:0] ? myVec_7 : _GEN_560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_562 = 7'h8 == _myNewVec_124_T_3[6:0] ? myVec_8 : _GEN_561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_563 = 7'h9 == _myNewVec_124_T_3[6:0] ? myVec_9 : _GEN_562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_564 = 7'ha == _myNewVec_124_T_3[6:0] ? myVec_10 : _GEN_563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_565 = 7'hb == _myNewVec_124_T_3[6:0] ? myVec_11 : _GEN_564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_566 = 7'hc == _myNewVec_124_T_3[6:0] ? myVec_12 : _GEN_565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_567 = 7'hd == _myNewVec_124_T_3[6:0] ? myVec_13 : _GEN_566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_568 = 7'he == _myNewVec_124_T_3[6:0] ? myVec_14 : _GEN_567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_569 = 7'hf == _myNewVec_124_T_3[6:0] ? myVec_15 : _GEN_568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_570 = 7'h10 == _myNewVec_124_T_3[6:0] ? myVec_16 : _GEN_569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_571 = 7'h11 == _myNewVec_124_T_3[6:0] ? myVec_17 : _GEN_570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_572 = 7'h12 == _myNewVec_124_T_3[6:0] ? myVec_18 : _GEN_571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_573 = 7'h13 == _myNewVec_124_T_3[6:0] ? myVec_19 : _GEN_572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_574 = 7'h14 == _myNewVec_124_T_3[6:0] ? myVec_20 : _GEN_573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_575 = 7'h15 == _myNewVec_124_T_3[6:0] ? myVec_21 : _GEN_574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_576 = 7'h16 == _myNewVec_124_T_3[6:0] ? myVec_22 : _GEN_575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_577 = 7'h17 == _myNewVec_124_T_3[6:0] ? myVec_23 : _GEN_576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_578 = 7'h18 == _myNewVec_124_T_3[6:0] ? myVec_24 : _GEN_577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_579 = 7'h19 == _myNewVec_124_T_3[6:0] ? myVec_25 : _GEN_578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_580 = 7'h1a == _myNewVec_124_T_3[6:0] ? myVec_26 : _GEN_579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_581 = 7'h1b == _myNewVec_124_T_3[6:0] ? myVec_27 : _GEN_580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_582 = 7'h1c == _myNewVec_124_T_3[6:0] ? myVec_28 : _GEN_581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_583 = 7'h1d == _myNewVec_124_T_3[6:0] ? myVec_29 : _GEN_582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_584 = 7'h1e == _myNewVec_124_T_3[6:0] ? myVec_30 : _GEN_583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_585 = 7'h1f == _myNewVec_124_T_3[6:0] ? myVec_31 : _GEN_584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_586 = 7'h20 == _myNewVec_124_T_3[6:0] ? myVec_32 : _GEN_585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_587 = 7'h21 == _myNewVec_124_T_3[6:0] ? myVec_33 : _GEN_586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_588 = 7'h22 == _myNewVec_124_T_3[6:0] ? myVec_34 : _GEN_587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_589 = 7'h23 == _myNewVec_124_T_3[6:0] ? myVec_35 : _GEN_588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_590 = 7'h24 == _myNewVec_124_T_3[6:0] ? myVec_36 : _GEN_589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_591 = 7'h25 == _myNewVec_124_T_3[6:0] ? myVec_37 : _GEN_590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_592 = 7'h26 == _myNewVec_124_T_3[6:0] ? myVec_38 : _GEN_591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_593 = 7'h27 == _myNewVec_124_T_3[6:0] ? myVec_39 : _GEN_592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_594 = 7'h28 == _myNewVec_124_T_3[6:0] ? myVec_40 : _GEN_593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_595 = 7'h29 == _myNewVec_124_T_3[6:0] ? myVec_41 : _GEN_594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_596 = 7'h2a == _myNewVec_124_T_3[6:0] ? myVec_42 : _GEN_595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_597 = 7'h2b == _myNewVec_124_T_3[6:0] ? myVec_43 : _GEN_596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_598 = 7'h2c == _myNewVec_124_T_3[6:0] ? myVec_44 : _GEN_597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_599 = 7'h2d == _myNewVec_124_T_3[6:0] ? myVec_45 : _GEN_598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_600 = 7'h2e == _myNewVec_124_T_3[6:0] ? myVec_46 : _GEN_599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_601 = 7'h2f == _myNewVec_124_T_3[6:0] ? myVec_47 : _GEN_600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_602 = 7'h30 == _myNewVec_124_T_3[6:0] ? myVec_48 : _GEN_601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_603 = 7'h31 == _myNewVec_124_T_3[6:0] ? myVec_49 : _GEN_602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_604 = 7'h32 == _myNewVec_124_T_3[6:0] ? myVec_50 : _GEN_603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_605 = 7'h33 == _myNewVec_124_T_3[6:0] ? myVec_51 : _GEN_604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_606 = 7'h34 == _myNewVec_124_T_3[6:0] ? myVec_52 : _GEN_605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_607 = 7'h35 == _myNewVec_124_T_3[6:0] ? myVec_53 : _GEN_606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_608 = 7'h36 == _myNewVec_124_T_3[6:0] ? myVec_54 : _GEN_607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_609 = 7'h37 == _myNewVec_124_T_3[6:0] ? myVec_55 : _GEN_608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_610 = 7'h38 == _myNewVec_124_T_3[6:0] ? myVec_56 : _GEN_609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_611 = 7'h39 == _myNewVec_124_T_3[6:0] ? myVec_57 : _GEN_610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_612 = 7'h3a == _myNewVec_124_T_3[6:0] ? myVec_58 : _GEN_611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_613 = 7'h3b == _myNewVec_124_T_3[6:0] ? myVec_59 : _GEN_612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_614 = 7'h3c == _myNewVec_124_T_3[6:0] ? myVec_60 : _GEN_613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_615 = 7'h3d == _myNewVec_124_T_3[6:0] ? myVec_61 : _GEN_614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_616 = 7'h3e == _myNewVec_124_T_3[6:0] ? myVec_62 : _GEN_615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_617 = 7'h3f == _myNewVec_124_T_3[6:0] ? myVec_63 : _GEN_616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_618 = 7'h40 == _myNewVec_124_T_3[6:0] ? myVec_64 : _GEN_617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_619 = 7'h41 == _myNewVec_124_T_3[6:0] ? myVec_65 : _GEN_618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_620 = 7'h42 == _myNewVec_124_T_3[6:0] ? myVec_66 : _GEN_619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_621 = 7'h43 == _myNewVec_124_T_3[6:0] ? myVec_67 : _GEN_620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_622 = 7'h44 == _myNewVec_124_T_3[6:0] ? myVec_68 : _GEN_621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_623 = 7'h45 == _myNewVec_124_T_3[6:0] ? myVec_69 : _GEN_622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_624 = 7'h46 == _myNewVec_124_T_3[6:0] ? myVec_70 : _GEN_623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_625 = 7'h47 == _myNewVec_124_T_3[6:0] ? myVec_71 : _GEN_624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_626 = 7'h48 == _myNewVec_124_T_3[6:0] ? myVec_72 : _GEN_625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_627 = 7'h49 == _myNewVec_124_T_3[6:0] ? myVec_73 : _GEN_626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_628 = 7'h4a == _myNewVec_124_T_3[6:0] ? myVec_74 : _GEN_627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_629 = 7'h4b == _myNewVec_124_T_3[6:0] ? myVec_75 : _GEN_628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_630 = 7'h4c == _myNewVec_124_T_3[6:0] ? myVec_76 : _GEN_629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_631 = 7'h4d == _myNewVec_124_T_3[6:0] ? myVec_77 : _GEN_630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_632 = 7'h4e == _myNewVec_124_T_3[6:0] ? myVec_78 : _GEN_631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_633 = 7'h4f == _myNewVec_124_T_3[6:0] ? myVec_79 : _GEN_632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_634 = 7'h50 == _myNewVec_124_T_3[6:0] ? myVec_80 : _GEN_633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_635 = 7'h51 == _myNewVec_124_T_3[6:0] ? myVec_81 : _GEN_634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_636 = 7'h52 == _myNewVec_124_T_3[6:0] ? myVec_82 : _GEN_635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_637 = 7'h53 == _myNewVec_124_T_3[6:0] ? myVec_83 : _GEN_636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_638 = 7'h54 == _myNewVec_124_T_3[6:0] ? myVec_84 : _GEN_637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_639 = 7'h55 == _myNewVec_124_T_3[6:0] ? myVec_85 : _GEN_638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_640 = 7'h56 == _myNewVec_124_T_3[6:0] ? myVec_86 : _GEN_639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_641 = 7'h57 == _myNewVec_124_T_3[6:0] ? myVec_87 : _GEN_640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_642 = 7'h58 == _myNewVec_124_T_3[6:0] ? myVec_88 : _GEN_641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_643 = 7'h59 == _myNewVec_124_T_3[6:0] ? myVec_89 : _GEN_642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_644 = 7'h5a == _myNewVec_124_T_3[6:0] ? myVec_90 : _GEN_643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_645 = 7'h5b == _myNewVec_124_T_3[6:0] ? myVec_91 : _GEN_644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_646 = 7'h5c == _myNewVec_124_T_3[6:0] ? myVec_92 : _GEN_645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_647 = 7'h5d == _myNewVec_124_T_3[6:0] ? myVec_93 : _GEN_646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_648 = 7'h5e == _myNewVec_124_T_3[6:0] ? myVec_94 : _GEN_647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_649 = 7'h5f == _myNewVec_124_T_3[6:0] ? myVec_95 : _GEN_648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_650 = 7'h60 == _myNewVec_124_T_3[6:0] ? myVec_96 : _GEN_649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_651 = 7'h61 == _myNewVec_124_T_3[6:0] ? myVec_97 : _GEN_650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_652 = 7'h62 == _myNewVec_124_T_3[6:0] ? myVec_98 : _GEN_651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_653 = 7'h63 == _myNewVec_124_T_3[6:0] ? myVec_99 : _GEN_652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_654 = 7'h64 == _myNewVec_124_T_3[6:0] ? myVec_100 : _GEN_653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_655 = 7'h65 == _myNewVec_124_T_3[6:0] ? myVec_101 : _GEN_654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_656 = 7'h66 == _myNewVec_124_T_3[6:0] ? myVec_102 : _GEN_655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_657 = 7'h67 == _myNewVec_124_T_3[6:0] ? myVec_103 : _GEN_656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_658 = 7'h68 == _myNewVec_124_T_3[6:0] ? myVec_104 : _GEN_657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_659 = 7'h69 == _myNewVec_124_T_3[6:0] ? myVec_105 : _GEN_658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_660 = 7'h6a == _myNewVec_124_T_3[6:0] ? myVec_106 : _GEN_659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_661 = 7'h6b == _myNewVec_124_T_3[6:0] ? myVec_107 : _GEN_660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_662 = 7'h6c == _myNewVec_124_T_3[6:0] ? myVec_108 : _GEN_661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_663 = 7'h6d == _myNewVec_124_T_3[6:0] ? myVec_109 : _GEN_662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_664 = 7'h6e == _myNewVec_124_T_3[6:0] ? myVec_110 : _GEN_663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_665 = 7'h6f == _myNewVec_124_T_3[6:0] ? myVec_111 : _GEN_664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_666 = 7'h70 == _myNewVec_124_T_3[6:0] ? myVec_112 : _GEN_665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_667 = 7'h71 == _myNewVec_124_T_3[6:0] ? myVec_113 : _GEN_666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_668 = 7'h72 == _myNewVec_124_T_3[6:0] ? myVec_114 : _GEN_667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_669 = 7'h73 == _myNewVec_124_T_3[6:0] ? myVec_115 : _GEN_668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_670 = 7'h74 == _myNewVec_124_T_3[6:0] ? myVec_116 : _GEN_669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_671 = 7'h75 == _myNewVec_124_T_3[6:0] ? myVec_117 : _GEN_670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_672 = 7'h76 == _myNewVec_124_T_3[6:0] ? myVec_118 : _GEN_671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_673 = 7'h77 == _myNewVec_124_T_3[6:0] ? myVec_119 : _GEN_672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_674 = 7'h78 == _myNewVec_124_T_3[6:0] ? myVec_120 : _GEN_673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_675 = 7'h79 == _myNewVec_124_T_3[6:0] ? myVec_121 : _GEN_674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_676 = 7'h7a == _myNewVec_124_T_3[6:0] ? myVec_122 : _GEN_675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_677 = 7'h7b == _myNewVec_124_T_3[6:0] ? myVec_123 : _GEN_676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_678 = 7'h7c == _myNewVec_124_T_3[6:0] ? myVec_124 : _GEN_677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_679 = 7'h7d == _myNewVec_124_T_3[6:0] ? myVec_125 : _GEN_678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_680 = 7'h7e == _myNewVec_124_T_3[6:0] ? myVec_126 : _GEN_679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_124 = 7'h7f == _myNewVec_124_T_3[6:0] ? myVec_127 : _GEN_680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_123_T_3 = _myNewVec_127_T_1 + 16'h4; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_683 = 7'h1 == _myNewVec_123_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_684 = 7'h2 == _myNewVec_123_T_3[6:0] ? myVec_2 : _GEN_683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_685 = 7'h3 == _myNewVec_123_T_3[6:0] ? myVec_3 : _GEN_684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_686 = 7'h4 == _myNewVec_123_T_3[6:0] ? myVec_4 : _GEN_685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_687 = 7'h5 == _myNewVec_123_T_3[6:0] ? myVec_5 : _GEN_686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_688 = 7'h6 == _myNewVec_123_T_3[6:0] ? myVec_6 : _GEN_687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_689 = 7'h7 == _myNewVec_123_T_3[6:0] ? myVec_7 : _GEN_688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_690 = 7'h8 == _myNewVec_123_T_3[6:0] ? myVec_8 : _GEN_689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_691 = 7'h9 == _myNewVec_123_T_3[6:0] ? myVec_9 : _GEN_690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_692 = 7'ha == _myNewVec_123_T_3[6:0] ? myVec_10 : _GEN_691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_693 = 7'hb == _myNewVec_123_T_3[6:0] ? myVec_11 : _GEN_692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_694 = 7'hc == _myNewVec_123_T_3[6:0] ? myVec_12 : _GEN_693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_695 = 7'hd == _myNewVec_123_T_3[6:0] ? myVec_13 : _GEN_694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_696 = 7'he == _myNewVec_123_T_3[6:0] ? myVec_14 : _GEN_695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_697 = 7'hf == _myNewVec_123_T_3[6:0] ? myVec_15 : _GEN_696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_698 = 7'h10 == _myNewVec_123_T_3[6:0] ? myVec_16 : _GEN_697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_699 = 7'h11 == _myNewVec_123_T_3[6:0] ? myVec_17 : _GEN_698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_700 = 7'h12 == _myNewVec_123_T_3[6:0] ? myVec_18 : _GEN_699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_701 = 7'h13 == _myNewVec_123_T_3[6:0] ? myVec_19 : _GEN_700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_702 = 7'h14 == _myNewVec_123_T_3[6:0] ? myVec_20 : _GEN_701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_703 = 7'h15 == _myNewVec_123_T_3[6:0] ? myVec_21 : _GEN_702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_704 = 7'h16 == _myNewVec_123_T_3[6:0] ? myVec_22 : _GEN_703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_705 = 7'h17 == _myNewVec_123_T_3[6:0] ? myVec_23 : _GEN_704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_706 = 7'h18 == _myNewVec_123_T_3[6:0] ? myVec_24 : _GEN_705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_707 = 7'h19 == _myNewVec_123_T_3[6:0] ? myVec_25 : _GEN_706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_708 = 7'h1a == _myNewVec_123_T_3[6:0] ? myVec_26 : _GEN_707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_709 = 7'h1b == _myNewVec_123_T_3[6:0] ? myVec_27 : _GEN_708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_710 = 7'h1c == _myNewVec_123_T_3[6:0] ? myVec_28 : _GEN_709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_711 = 7'h1d == _myNewVec_123_T_3[6:0] ? myVec_29 : _GEN_710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_712 = 7'h1e == _myNewVec_123_T_3[6:0] ? myVec_30 : _GEN_711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_713 = 7'h1f == _myNewVec_123_T_3[6:0] ? myVec_31 : _GEN_712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_714 = 7'h20 == _myNewVec_123_T_3[6:0] ? myVec_32 : _GEN_713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_715 = 7'h21 == _myNewVec_123_T_3[6:0] ? myVec_33 : _GEN_714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_716 = 7'h22 == _myNewVec_123_T_3[6:0] ? myVec_34 : _GEN_715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_717 = 7'h23 == _myNewVec_123_T_3[6:0] ? myVec_35 : _GEN_716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_718 = 7'h24 == _myNewVec_123_T_3[6:0] ? myVec_36 : _GEN_717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_719 = 7'h25 == _myNewVec_123_T_3[6:0] ? myVec_37 : _GEN_718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_720 = 7'h26 == _myNewVec_123_T_3[6:0] ? myVec_38 : _GEN_719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_721 = 7'h27 == _myNewVec_123_T_3[6:0] ? myVec_39 : _GEN_720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_722 = 7'h28 == _myNewVec_123_T_3[6:0] ? myVec_40 : _GEN_721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_723 = 7'h29 == _myNewVec_123_T_3[6:0] ? myVec_41 : _GEN_722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_724 = 7'h2a == _myNewVec_123_T_3[6:0] ? myVec_42 : _GEN_723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_725 = 7'h2b == _myNewVec_123_T_3[6:0] ? myVec_43 : _GEN_724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_726 = 7'h2c == _myNewVec_123_T_3[6:0] ? myVec_44 : _GEN_725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_727 = 7'h2d == _myNewVec_123_T_3[6:0] ? myVec_45 : _GEN_726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_728 = 7'h2e == _myNewVec_123_T_3[6:0] ? myVec_46 : _GEN_727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_729 = 7'h2f == _myNewVec_123_T_3[6:0] ? myVec_47 : _GEN_728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_730 = 7'h30 == _myNewVec_123_T_3[6:0] ? myVec_48 : _GEN_729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_731 = 7'h31 == _myNewVec_123_T_3[6:0] ? myVec_49 : _GEN_730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_732 = 7'h32 == _myNewVec_123_T_3[6:0] ? myVec_50 : _GEN_731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_733 = 7'h33 == _myNewVec_123_T_3[6:0] ? myVec_51 : _GEN_732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_734 = 7'h34 == _myNewVec_123_T_3[6:0] ? myVec_52 : _GEN_733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_735 = 7'h35 == _myNewVec_123_T_3[6:0] ? myVec_53 : _GEN_734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_736 = 7'h36 == _myNewVec_123_T_3[6:0] ? myVec_54 : _GEN_735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_737 = 7'h37 == _myNewVec_123_T_3[6:0] ? myVec_55 : _GEN_736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_738 = 7'h38 == _myNewVec_123_T_3[6:0] ? myVec_56 : _GEN_737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_739 = 7'h39 == _myNewVec_123_T_3[6:0] ? myVec_57 : _GEN_738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_740 = 7'h3a == _myNewVec_123_T_3[6:0] ? myVec_58 : _GEN_739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_741 = 7'h3b == _myNewVec_123_T_3[6:0] ? myVec_59 : _GEN_740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_742 = 7'h3c == _myNewVec_123_T_3[6:0] ? myVec_60 : _GEN_741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_743 = 7'h3d == _myNewVec_123_T_3[6:0] ? myVec_61 : _GEN_742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_744 = 7'h3e == _myNewVec_123_T_3[6:0] ? myVec_62 : _GEN_743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_745 = 7'h3f == _myNewVec_123_T_3[6:0] ? myVec_63 : _GEN_744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_746 = 7'h40 == _myNewVec_123_T_3[6:0] ? myVec_64 : _GEN_745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_747 = 7'h41 == _myNewVec_123_T_3[6:0] ? myVec_65 : _GEN_746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_748 = 7'h42 == _myNewVec_123_T_3[6:0] ? myVec_66 : _GEN_747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_749 = 7'h43 == _myNewVec_123_T_3[6:0] ? myVec_67 : _GEN_748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_750 = 7'h44 == _myNewVec_123_T_3[6:0] ? myVec_68 : _GEN_749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_751 = 7'h45 == _myNewVec_123_T_3[6:0] ? myVec_69 : _GEN_750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_752 = 7'h46 == _myNewVec_123_T_3[6:0] ? myVec_70 : _GEN_751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_753 = 7'h47 == _myNewVec_123_T_3[6:0] ? myVec_71 : _GEN_752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_754 = 7'h48 == _myNewVec_123_T_3[6:0] ? myVec_72 : _GEN_753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_755 = 7'h49 == _myNewVec_123_T_3[6:0] ? myVec_73 : _GEN_754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_756 = 7'h4a == _myNewVec_123_T_3[6:0] ? myVec_74 : _GEN_755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_757 = 7'h4b == _myNewVec_123_T_3[6:0] ? myVec_75 : _GEN_756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_758 = 7'h4c == _myNewVec_123_T_3[6:0] ? myVec_76 : _GEN_757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_759 = 7'h4d == _myNewVec_123_T_3[6:0] ? myVec_77 : _GEN_758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_760 = 7'h4e == _myNewVec_123_T_3[6:0] ? myVec_78 : _GEN_759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_761 = 7'h4f == _myNewVec_123_T_3[6:0] ? myVec_79 : _GEN_760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_762 = 7'h50 == _myNewVec_123_T_3[6:0] ? myVec_80 : _GEN_761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_763 = 7'h51 == _myNewVec_123_T_3[6:0] ? myVec_81 : _GEN_762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_764 = 7'h52 == _myNewVec_123_T_3[6:0] ? myVec_82 : _GEN_763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_765 = 7'h53 == _myNewVec_123_T_3[6:0] ? myVec_83 : _GEN_764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_766 = 7'h54 == _myNewVec_123_T_3[6:0] ? myVec_84 : _GEN_765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_767 = 7'h55 == _myNewVec_123_T_3[6:0] ? myVec_85 : _GEN_766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_768 = 7'h56 == _myNewVec_123_T_3[6:0] ? myVec_86 : _GEN_767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_769 = 7'h57 == _myNewVec_123_T_3[6:0] ? myVec_87 : _GEN_768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_770 = 7'h58 == _myNewVec_123_T_3[6:0] ? myVec_88 : _GEN_769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_771 = 7'h59 == _myNewVec_123_T_3[6:0] ? myVec_89 : _GEN_770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_772 = 7'h5a == _myNewVec_123_T_3[6:0] ? myVec_90 : _GEN_771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_773 = 7'h5b == _myNewVec_123_T_3[6:0] ? myVec_91 : _GEN_772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_774 = 7'h5c == _myNewVec_123_T_3[6:0] ? myVec_92 : _GEN_773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_775 = 7'h5d == _myNewVec_123_T_3[6:0] ? myVec_93 : _GEN_774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_776 = 7'h5e == _myNewVec_123_T_3[6:0] ? myVec_94 : _GEN_775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_777 = 7'h5f == _myNewVec_123_T_3[6:0] ? myVec_95 : _GEN_776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_778 = 7'h60 == _myNewVec_123_T_3[6:0] ? myVec_96 : _GEN_777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_779 = 7'h61 == _myNewVec_123_T_3[6:0] ? myVec_97 : _GEN_778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_780 = 7'h62 == _myNewVec_123_T_3[6:0] ? myVec_98 : _GEN_779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_781 = 7'h63 == _myNewVec_123_T_3[6:0] ? myVec_99 : _GEN_780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_782 = 7'h64 == _myNewVec_123_T_3[6:0] ? myVec_100 : _GEN_781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_783 = 7'h65 == _myNewVec_123_T_3[6:0] ? myVec_101 : _GEN_782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_784 = 7'h66 == _myNewVec_123_T_3[6:0] ? myVec_102 : _GEN_783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_785 = 7'h67 == _myNewVec_123_T_3[6:0] ? myVec_103 : _GEN_784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_786 = 7'h68 == _myNewVec_123_T_3[6:0] ? myVec_104 : _GEN_785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_787 = 7'h69 == _myNewVec_123_T_3[6:0] ? myVec_105 : _GEN_786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_788 = 7'h6a == _myNewVec_123_T_3[6:0] ? myVec_106 : _GEN_787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_789 = 7'h6b == _myNewVec_123_T_3[6:0] ? myVec_107 : _GEN_788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_790 = 7'h6c == _myNewVec_123_T_3[6:0] ? myVec_108 : _GEN_789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_791 = 7'h6d == _myNewVec_123_T_3[6:0] ? myVec_109 : _GEN_790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_792 = 7'h6e == _myNewVec_123_T_3[6:0] ? myVec_110 : _GEN_791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_793 = 7'h6f == _myNewVec_123_T_3[6:0] ? myVec_111 : _GEN_792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_794 = 7'h70 == _myNewVec_123_T_3[6:0] ? myVec_112 : _GEN_793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_795 = 7'h71 == _myNewVec_123_T_3[6:0] ? myVec_113 : _GEN_794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_796 = 7'h72 == _myNewVec_123_T_3[6:0] ? myVec_114 : _GEN_795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_797 = 7'h73 == _myNewVec_123_T_3[6:0] ? myVec_115 : _GEN_796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_798 = 7'h74 == _myNewVec_123_T_3[6:0] ? myVec_116 : _GEN_797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_799 = 7'h75 == _myNewVec_123_T_3[6:0] ? myVec_117 : _GEN_798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_800 = 7'h76 == _myNewVec_123_T_3[6:0] ? myVec_118 : _GEN_799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_801 = 7'h77 == _myNewVec_123_T_3[6:0] ? myVec_119 : _GEN_800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_802 = 7'h78 == _myNewVec_123_T_3[6:0] ? myVec_120 : _GEN_801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_803 = 7'h79 == _myNewVec_123_T_3[6:0] ? myVec_121 : _GEN_802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_804 = 7'h7a == _myNewVec_123_T_3[6:0] ? myVec_122 : _GEN_803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_805 = 7'h7b == _myNewVec_123_T_3[6:0] ? myVec_123 : _GEN_804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_806 = 7'h7c == _myNewVec_123_T_3[6:0] ? myVec_124 : _GEN_805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_807 = 7'h7d == _myNewVec_123_T_3[6:0] ? myVec_125 : _GEN_806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_808 = 7'h7e == _myNewVec_123_T_3[6:0] ? myVec_126 : _GEN_807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_123 = 7'h7f == _myNewVec_123_T_3[6:0] ? myVec_127 : _GEN_808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_122_T_3 = _myNewVec_127_T_1 + 16'h5; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_811 = 7'h1 == _myNewVec_122_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_812 = 7'h2 == _myNewVec_122_T_3[6:0] ? myVec_2 : _GEN_811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_813 = 7'h3 == _myNewVec_122_T_3[6:0] ? myVec_3 : _GEN_812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_814 = 7'h4 == _myNewVec_122_T_3[6:0] ? myVec_4 : _GEN_813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_815 = 7'h5 == _myNewVec_122_T_3[6:0] ? myVec_5 : _GEN_814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_816 = 7'h6 == _myNewVec_122_T_3[6:0] ? myVec_6 : _GEN_815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_817 = 7'h7 == _myNewVec_122_T_3[6:0] ? myVec_7 : _GEN_816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_818 = 7'h8 == _myNewVec_122_T_3[6:0] ? myVec_8 : _GEN_817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_819 = 7'h9 == _myNewVec_122_T_3[6:0] ? myVec_9 : _GEN_818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_820 = 7'ha == _myNewVec_122_T_3[6:0] ? myVec_10 : _GEN_819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_821 = 7'hb == _myNewVec_122_T_3[6:0] ? myVec_11 : _GEN_820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_822 = 7'hc == _myNewVec_122_T_3[6:0] ? myVec_12 : _GEN_821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_823 = 7'hd == _myNewVec_122_T_3[6:0] ? myVec_13 : _GEN_822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_824 = 7'he == _myNewVec_122_T_3[6:0] ? myVec_14 : _GEN_823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_825 = 7'hf == _myNewVec_122_T_3[6:0] ? myVec_15 : _GEN_824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_826 = 7'h10 == _myNewVec_122_T_3[6:0] ? myVec_16 : _GEN_825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_827 = 7'h11 == _myNewVec_122_T_3[6:0] ? myVec_17 : _GEN_826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_828 = 7'h12 == _myNewVec_122_T_3[6:0] ? myVec_18 : _GEN_827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_829 = 7'h13 == _myNewVec_122_T_3[6:0] ? myVec_19 : _GEN_828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_830 = 7'h14 == _myNewVec_122_T_3[6:0] ? myVec_20 : _GEN_829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_831 = 7'h15 == _myNewVec_122_T_3[6:0] ? myVec_21 : _GEN_830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_832 = 7'h16 == _myNewVec_122_T_3[6:0] ? myVec_22 : _GEN_831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_833 = 7'h17 == _myNewVec_122_T_3[6:0] ? myVec_23 : _GEN_832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_834 = 7'h18 == _myNewVec_122_T_3[6:0] ? myVec_24 : _GEN_833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_835 = 7'h19 == _myNewVec_122_T_3[6:0] ? myVec_25 : _GEN_834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_836 = 7'h1a == _myNewVec_122_T_3[6:0] ? myVec_26 : _GEN_835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_837 = 7'h1b == _myNewVec_122_T_3[6:0] ? myVec_27 : _GEN_836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_838 = 7'h1c == _myNewVec_122_T_3[6:0] ? myVec_28 : _GEN_837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_839 = 7'h1d == _myNewVec_122_T_3[6:0] ? myVec_29 : _GEN_838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_840 = 7'h1e == _myNewVec_122_T_3[6:0] ? myVec_30 : _GEN_839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_841 = 7'h1f == _myNewVec_122_T_3[6:0] ? myVec_31 : _GEN_840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_842 = 7'h20 == _myNewVec_122_T_3[6:0] ? myVec_32 : _GEN_841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_843 = 7'h21 == _myNewVec_122_T_3[6:0] ? myVec_33 : _GEN_842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_844 = 7'h22 == _myNewVec_122_T_3[6:0] ? myVec_34 : _GEN_843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_845 = 7'h23 == _myNewVec_122_T_3[6:0] ? myVec_35 : _GEN_844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_846 = 7'h24 == _myNewVec_122_T_3[6:0] ? myVec_36 : _GEN_845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_847 = 7'h25 == _myNewVec_122_T_3[6:0] ? myVec_37 : _GEN_846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_848 = 7'h26 == _myNewVec_122_T_3[6:0] ? myVec_38 : _GEN_847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_849 = 7'h27 == _myNewVec_122_T_3[6:0] ? myVec_39 : _GEN_848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_850 = 7'h28 == _myNewVec_122_T_3[6:0] ? myVec_40 : _GEN_849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_851 = 7'h29 == _myNewVec_122_T_3[6:0] ? myVec_41 : _GEN_850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_852 = 7'h2a == _myNewVec_122_T_3[6:0] ? myVec_42 : _GEN_851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_853 = 7'h2b == _myNewVec_122_T_3[6:0] ? myVec_43 : _GEN_852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_854 = 7'h2c == _myNewVec_122_T_3[6:0] ? myVec_44 : _GEN_853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_855 = 7'h2d == _myNewVec_122_T_3[6:0] ? myVec_45 : _GEN_854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_856 = 7'h2e == _myNewVec_122_T_3[6:0] ? myVec_46 : _GEN_855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_857 = 7'h2f == _myNewVec_122_T_3[6:0] ? myVec_47 : _GEN_856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_858 = 7'h30 == _myNewVec_122_T_3[6:0] ? myVec_48 : _GEN_857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_859 = 7'h31 == _myNewVec_122_T_3[6:0] ? myVec_49 : _GEN_858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_860 = 7'h32 == _myNewVec_122_T_3[6:0] ? myVec_50 : _GEN_859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_861 = 7'h33 == _myNewVec_122_T_3[6:0] ? myVec_51 : _GEN_860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_862 = 7'h34 == _myNewVec_122_T_3[6:0] ? myVec_52 : _GEN_861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_863 = 7'h35 == _myNewVec_122_T_3[6:0] ? myVec_53 : _GEN_862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_864 = 7'h36 == _myNewVec_122_T_3[6:0] ? myVec_54 : _GEN_863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_865 = 7'h37 == _myNewVec_122_T_3[6:0] ? myVec_55 : _GEN_864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_866 = 7'h38 == _myNewVec_122_T_3[6:0] ? myVec_56 : _GEN_865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_867 = 7'h39 == _myNewVec_122_T_3[6:0] ? myVec_57 : _GEN_866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_868 = 7'h3a == _myNewVec_122_T_3[6:0] ? myVec_58 : _GEN_867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_869 = 7'h3b == _myNewVec_122_T_3[6:0] ? myVec_59 : _GEN_868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_870 = 7'h3c == _myNewVec_122_T_3[6:0] ? myVec_60 : _GEN_869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_871 = 7'h3d == _myNewVec_122_T_3[6:0] ? myVec_61 : _GEN_870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_872 = 7'h3e == _myNewVec_122_T_3[6:0] ? myVec_62 : _GEN_871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_873 = 7'h3f == _myNewVec_122_T_3[6:0] ? myVec_63 : _GEN_872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_874 = 7'h40 == _myNewVec_122_T_3[6:0] ? myVec_64 : _GEN_873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_875 = 7'h41 == _myNewVec_122_T_3[6:0] ? myVec_65 : _GEN_874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_876 = 7'h42 == _myNewVec_122_T_3[6:0] ? myVec_66 : _GEN_875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_877 = 7'h43 == _myNewVec_122_T_3[6:0] ? myVec_67 : _GEN_876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_878 = 7'h44 == _myNewVec_122_T_3[6:0] ? myVec_68 : _GEN_877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_879 = 7'h45 == _myNewVec_122_T_3[6:0] ? myVec_69 : _GEN_878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_880 = 7'h46 == _myNewVec_122_T_3[6:0] ? myVec_70 : _GEN_879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_881 = 7'h47 == _myNewVec_122_T_3[6:0] ? myVec_71 : _GEN_880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_882 = 7'h48 == _myNewVec_122_T_3[6:0] ? myVec_72 : _GEN_881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_883 = 7'h49 == _myNewVec_122_T_3[6:0] ? myVec_73 : _GEN_882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_884 = 7'h4a == _myNewVec_122_T_3[6:0] ? myVec_74 : _GEN_883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_885 = 7'h4b == _myNewVec_122_T_3[6:0] ? myVec_75 : _GEN_884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_886 = 7'h4c == _myNewVec_122_T_3[6:0] ? myVec_76 : _GEN_885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_887 = 7'h4d == _myNewVec_122_T_3[6:0] ? myVec_77 : _GEN_886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_888 = 7'h4e == _myNewVec_122_T_3[6:0] ? myVec_78 : _GEN_887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_889 = 7'h4f == _myNewVec_122_T_3[6:0] ? myVec_79 : _GEN_888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_890 = 7'h50 == _myNewVec_122_T_3[6:0] ? myVec_80 : _GEN_889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_891 = 7'h51 == _myNewVec_122_T_3[6:0] ? myVec_81 : _GEN_890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_892 = 7'h52 == _myNewVec_122_T_3[6:0] ? myVec_82 : _GEN_891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_893 = 7'h53 == _myNewVec_122_T_3[6:0] ? myVec_83 : _GEN_892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_894 = 7'h54 == _myNewVec_122_T_3[6:0] ? myVec_84 : _GEN_893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_895 = 7'h55 == _myNewVec_122_T_3[6:0] ? myVec_85 : _GEN_894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_896 = 7'h56 == _myNewVec_122_T_3[6:0] ? myVec_86 : _GEN_895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_897 = 7'h57 == _myNewVec_122_T_3[6:0] ? myVec_87 : _GEN_896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_898 = 7'h58 == _myNewVec_122_T_3[6:0] ? myVec_88 : _GEN_897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_899 = 7'h59 == _myNewVec_122_T_3[6:0] ? myVec_89 : _GEN_898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_900 = 7'h5a == _myNewVec_122_T_3[6:0] ? myVec_90 : _GEN_899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_901 = 7'h5b == _myNewVec_122_T_3[6:0] ? myVec_91 : _GEN_900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_902 = 7'h5c == _myNewVec_122_T_3[6:0] ? myVec_92 : _GEN_901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_903 = 7'h5d == _myNewVec_122_T_3[6:0] ? myVec_93 : _GEN_902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_904 = 7'h5e == _myNewVec_122_T_3[6:0] ? myVec_94 : _GEN_903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_905 = 7'h5f == _myNewVec_122_T_3[6:0] ? myVec_95 : _GEN_904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_906 = 7'h60 == _myNewVec_122_T_3[6:0] ? myVec_96 : _GEN_905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_907 = 7'h61 == _myNewVec_122_T_3[6:0] ? myVec_97 : _GEN_906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_908 = 7'h62 == _myNewVec_122_T_3[6:0] ? myVec_98 : _GEN_907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_909 = 7'h63 == _myNewVec_122_T_3[6:0] ? myVec_99 : _GEN_908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_910 = 7'h64 == _myNewVec_122_T_3[6:0] ? myVec_100 : _GEN_909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_911 = 7'h65 == _myNewVec_122_T_3[6:0] ? myVec_101 : _GEN_910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_912 = 7'h66 == _myNewVec_122_T_3[6:0] ? myVec_102 : _GEN_911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_913 = 7'h67 == _myNewVec_122_T_3[6:0] ? myVec_103 : _GEN_912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_914 = 7'h68 == _myNewVec_122_T_3[6:0] ? myVec_104 : _GEN_913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_915 = 7'h69 == _myNewVec_122_T_3[6:0] ? myVec_105 : _GEN_914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_916 = 7'h6a == _myNewVec_122_T_3[6:0] ? myVec_106 : _GEN_915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_917 = 7'h6b == _myNewVec_122_T_3[6:0] ? myVec_107 : _GEN_916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_918 = 7'h6c == _myNewVec_122_T_3[6:0] ? myVec_108 : _GEN_917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_919 = 7'h6d == _myNewVec_122_T_3[6:0] ? myVec_109 : _GEN_918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_920 = 7'h6e == _myNewVec_122_T_3[6:0] ? myVec_110 : _GEN_919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_921 = 7'h6f == _myNewVec_122_T_3[6:0] ? myVec_111 : _GEN_920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_922 = 7'h70 == _myNewVec_122_T_3[6:0] ? myVec_112 : _GEN_921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_923 = 7'h71 == _myNewVec_122_T_3[6:0] ? myVec_113 : _GEN_922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_924 = 7'h72 == _myNewVec_122_T_3[6:0] ? myVec_114 : _GEN_923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_925 = 7'h73 == _myNewVec_122_T_3[6:0] ? myVec_115 : _GEN_924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_926 = 7'h74 == _myNewVec_122_T_3[6:0] ? myVec_116 : _GEN_925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_927 = 7'h75 == _myNewVec_122_T_3[6:0] ? myVec_117 : _GEN_926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_928 = 7'h76 == _myNewVec_122_T_3[6:0] ? myVec_118 : _GEN_927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_929 = 7'h77 == _myNewVec_122_T_3[6:0] ? myVec_119 : _GEN_928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_930 = 7'h78 == _myNewVec_122_T_3[6:0] ? myVec_120 : _GEN_929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_931 = 7'h79 == _myNewVec_122_T_3[6:0] ? myVec_121 : _GEN_930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_932 = 7'h7a == _myNewVec_122_T_3[6:0] ? myVec_122 : _GEN_931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_933 = 7'h7b == _myNewVec_122_T_3[6:0] ? myVec_123 : _GEN_932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_934 = 7'h7c == _myNewVec_122_T_3[6:0] ? myVec_124 : _GEN_933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_935 = 7'h7d == _myNewVec_122_T_3[6:0] ? myVec_125 : _GEN_934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_936 = 7'h7e == _myNewVec_122_T_3[6:0] ? myVec_126 : _GEN_935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_122 = 7'h7f == _myNewVec_122_T_3[6:0] ? myVec_127 : _GEN_936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_121_T_3 = _myNewVec_127_T_1 + 16'h6; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_939 = 7'h1 == _myNewVec_121_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_940 = 7'h2 == _myNewVec_121_T_3[6:0] ? myVec_2 : _GEN_939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_941 = 7'h3 == _myNewVec_121_T_3[6:0] ? myVec_3 : _GEN_940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_942 = 7'h4 == _myNewVec_121_T_3[6:0] ? myVec_4 : _GEN_941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_943 = 7'h5 == _myNewVec_121_T_3[6:0] ? myVec_5 : _GEN_942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_944 = 7'h6 == _myNewVec_121_T_3[6:0] ? myVec_6 : _GEN_943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_945 = 7'h7 == _myNewVec_121_T_3[6:0] ? myVec_7 : _GEN_944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_946 = 7'h8 == _myNewVec_121_T_3[6:0] ? myVec_8 : _GEN_945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_947 = 7'h9 == _myNewVec_121_T_3[6:0] ? myVec_9 : _GEN_946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_948 = 7'ha == _myNewVec_121_T_3[6:0] ? myVec_10 : _GEN_947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_949 = 7'hb == _myNewVec_121_T_3[6:0] ? myVec_11 : _GEN_948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_950 = 7'hc == _myNewVec_121_T_3[6:0] ? myVec_12 : _GEN_949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_951 = 7'hd == _myNewVec_121_T_3[6:0] ? myVec_13 : _GEN_950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_952 = 7'he == _myNewVec_121_T_3[6:0] ? myVec_14 : _GEN_951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_953 = 7'hf == _myNewVec_121_T_3[6:0] ? myVec_15 : _GEN_952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_954 = 7'h10 == _myNewVec_121_T_3[6:0] ? myVec_16 : _GEN_953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_955 = 7'h11 == _myNewVec_121_T_3[6:0] ? myVec_17 : _GEN_954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_956 = 7'h12 == _myNewVec_121_T_3[6:0] ? myVec_18 : _GEN_955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_957 = 7'h13 == _myNewVec_121_T_3[6:0] ? myVec_19 : _GEN_956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_958 = 7'h14 == _myNewVec_121_T_3[6:0] ? myVec_20 : _GEN_957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_959 = 7'h15 == _myNewVec_121_T_3[6:0] ? myVec_21 : _GEN_958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_960 = 7'h16 == _myNewVec_121_T_3[6:0] ? myVec_22 : _GEN_959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_961 = 7'h17 == _myNewVec_121_T_3[6:0] ? myVec_23 : _GEN_960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_962 = 7'h18 == _myNewVec_121_T_3[6:0] ? myVec_24 : _GEN_961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_963 = 7'h19 == _myNewVec_121_T_3[6:0] ? myVec_25 : _GEN_962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_964 = 7'h1a == _myNewVec_121_T_3[6:0] ? myVec_26 : _GEN_963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_965 = 7'h1b == _myNewVec_121_T_3[6:0] ? myVec_27 : _GEN_964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_966 = 7'h1c == _myNewVec_121_T_3[6:0] ? myVec_28 : _GEN_965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_967 = 7'h1d == _myNewVec_121_T_3[6:0] ? myVec_29 : _GEN_966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_968 = 7'h1e == _myNewVec_121_T_3[6:0] ? myVec_30 : _GEN_967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_969 = 7'h1f == _myNewVec_121_T_3[6:0] ? myVec_31 : _GEN_968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_970 = 7'h20 == _myNewVec_121_T_3[6:0] ? myVec_32 : _GEN_969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_971 = 7'h21 == _myNewVec_121_T_3[6:0] ? myVec_33 : _GEN_970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_972 = 7'h22 == _myNewVec_121_T_3[6:0] ? myVec_34 : _GEN_971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_973 = 7'h23 == _myNewVec_121_T_3[6:0] ? myVec_35 : _GEN_972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_974 = 7'h24 == _myNewVec_121_T_3[6:0] ? myVec_36 : _GEN_973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_975 = 7'h25 == _myNewVec_121_T_3[6:0] ? myVec_37 : _GEN_974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_976 = 7'h26 == _myNewVec_121_T_3[6:0] ? myVec_38 : _GEN_975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_977 = 7'h27 == _myNewVec_121_T_3[6:0] ? myVec_39 : _GEN_976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_978 = 7'h28 == _myNewVec_121_T_3[6:0] ? myVec_40 : _GEN_977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_979 = 7'h29 == _myNewVec_121_T_3[6:0] ? myVec_41 : _GEN_978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_980 = 7'h2a == _myNewVec_121_T_3[6:0] ? myVec_42 : _GEN_979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_981 = 7'h2b == _myNewVec_121_T_3[6:0] ? myVec_43 : _GEN_980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_982 = 7'h2c == _myNewVec_121_T_3[6:0] ? myVec_44 : _GEN_981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_983 = 7'h2d == _myNewVec_121_T_3[6:0] ? myVec_45 : _GEN_982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_984 = 7'h2e == _myNewVec_121_T_3[6:0] ? myVec_46 : _GEN_983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_985 = 7'h2f == _myNewVec_121_T_3[6:0] ? myVec_47 : _GEN_984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_986 = 7'h30 == _myNewVec_121_T_3[6:0] ? myVec_48 : _GEN_985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_987 = 7'h31 == _myNewVec_121_T_3[6:0] ? myVec_49 : _GEN_986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_988 = 7'h32 == _myNewVec_121_T_3[6:0] ? myVec_50 : _GEN_987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_989 = 7'h33 == _myNewVec_121_T_3[6:0] ? myVec_51 : _GEN_988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_990 = 7'h34 == _myNewVec_121_T_3[6:0] ? myVec_52 : _GEN_989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_991 = 7'h35 == _myNewVec_121_T_3[6:0] ? myVec_53 : _GEN_990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_992 = 7'h36 == _myNewVec_121_T_3[6:0] ? myVec_54 : _GEN_991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_993 = 7'h37 == _myNewVec_121_T_3[6:0] ? myVec_55 : _GEN_992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_994 = 7'h38 == _myNewVec_121_T_3[6:0] ? myVec_56 : _GEN_993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_995 = 7'h39 == _myNewVec_121_T_3[6:0] ? myVec_57 : _GEN_994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_996 = 7'h3a == _myNewVec_121_T_3[6:0] ? myVec_58 : _GEN_995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_997 = 7'h3b == _myNewVec_121_T_3[6:0] ? myVec_59 : _GEN_996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_998 = 7'h3c == _myNewVec_121_T_3[6:0] ? myVec_60 : _GEN_997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_999 = 7'h3d == _myNewVec_121_T_3[6:0] ? myVec_61 : _GEN_998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1000 = 7'h3e == _myNewVec_121_T_3[6:0] ? myVec_62 : _GEN_999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1001 = 7'h3f == _myNewVec_121_T_3[6:0] ? myVec_63 : _GEN_1000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1002 = 7'h40 == _myNewVec_121_T_3[6:0] ? myVec_64 : _GEN_1001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1003 = 7'h41 == _myNewVec_121_T_3[6:0] ? myVec_65 : _GEN_1002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1004 = 7'h42 == _myNewVec_121_T_3[6:0] ? myVec_66 : _GEN_1003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1005 = 7'h43 == _myNewVec_121_T_3[6:0] ? myVec_67 : _GEN_1004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1006 = 7'h44 == _myNewVec_121_T_3[6:0] ? myVec_68 : _GEN_1005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1007 = 7'h45 == _myNewVec_121_T_3[6:0] ? myVec_69 : _GEN_1006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1008 = 7'h46 == _myNewVec_121_T_3[6:0] ? myVec_70 : _GEN_1007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1009 = 7'h47 == _myNewVec_121_T_3[6:0] ? myVec_71 : _GEN_1008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1010 = 7'h48 == _myNewVec_121_T_3[6:0] ? myVec_72 : _GEN_1009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1011 = 7'h49 == _myNewVec_121_T_3[6:0] ? myVec_73 : _GEN_1010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1012 = 7'h4a == _myNewVec_121_T_3[6:0] ? myVec_74 : _GEN_1011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1013 = 7'h4b == _myNewVec_121_T_3[6:0] ? myVec_75 : _GEN_1012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1014 = 7'h4c == _myNewVec_121_T_3[6:0] ? myVec_76 : _GEN_1013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1015 = 7'h4d == _myNewVec_121_T_3[6:0] ? myVec_77 : _GEN_1014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1016 = 7'h4e == _myNewVec_121_T_3[6:0] ? myVec_78 : _GEN_1015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1017 = 7'h4f == _myNewVec_121_T_3[6:0] ? myVec_79 : _GEN_1016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1018 = 7'h50 == _myNewVec_121_T_3[6:0] ? myVec_80 : _GEN_1017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1019 = 7'h51 == _myNewVec_121_T_3[6:0] ? myVec_81 : _GEN_1018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1020 = 7'h52 == _myNewVec_121_T_3[6:0] ? myVec_82 : _GEN_1019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1021 = 7'h53 == _myNewVec_121_T_3[6:0] ? myVec_83 : _GEN_1020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1022 = 7'h54 == _myNewVec_121_T_3[6:0] ? myVec_84 : _GEN_1021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1023 = 7'h55 == _myNewVec_121_T_3[6:0] ? myVec_85 : _GEN_1022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1024 = 7'h56 == _myNewVec_121_T_3[6:0] ? myVec_86 : _GEN_1023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1025 = 7'h57 == _myNewVec_121_T_3[6:0] ? myVec_87 : _GEN_1024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1026 = 7'h58 == _myNewVec_121_T_3[6:0] ? myVec_88 : _GEN_1025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1027 = 7'h59 == _myNewVec_121_T_3[6:0] ? myVec_89 : _GEN_1026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1028 = 7'h5a == _myNewVec_121_T_3[6:0] ? myVec_90 : _GEN_1027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1029 = 7'h5b == _myNewVec_121_T_3[6:0] ? myVec_91 : _GEN_1028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1030 = 7'h5c == _myNewVec_121_T_3[6:0] ? myVec_92 : _GEN_1029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1031 = 7'h5d == _myNewVec_121_T_3[6:0] ? myVec_93 : _GEN_1030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1032 = 7'h5e == _myNewVec_121_T_3[6:0] ? myVec_94 : _GEN_1031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1033 = 7'h5f == _myNewVec_121_T_3[6:0] ? myVec_95 : _GEN_1032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1034 = 7'h60 == _myNewVec_121_T_3[6:0] ? myVec_96 : _GEN_1033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1035 = 7'h61 == _myNewVec_121_T_3[6:0] ? myVec_97 : _GEN_1034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1036 = 7'h62 == _myNewVec_121_T_3[6:0] ? myVec_98 : _GEN_1035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1037 = 7'h63 == _myNewVec_121_T_3[6:0] ? myVec_99 : _GEN_1036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1038 = 7'h64 == _myNewVec_121_T_3[6:0] ? myVec_100 : _GEN_1037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1039 = 7'h65 == _myNewVec_121_T_3[6:0] ? myVec_101 : _GEN_1038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1040 = 7'h66 == _myNewVec_121_T_3[6:0] ? myVec_102 : _GEN_1039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1041 = 7'h67 == _myNewVec_121_T_3[6:0] ? myVec_103 : _GEN_1040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1042 = 7'h68 == _myNewVec_121_T_3[6:0] ? myVec_104 : _GEN_1041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1043 = 7'h69 == _myNewVec_121_T_3[6:0] ? myVec_105 : _GEN_1042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1044 = 7'h6a == _myNewVec_121_T_3[6:0] ? myVec_106 : _GEN_1043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1045 = 7'h6b == _myNewVec_121_T_3[6:0] ? myVec_107 : _GEN_1044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1046 = 7'h6c == _myNewVec_121_T_3[6:0] ? myVec_108 : _GEN_1045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1047 = 7'h6d == _myNewVec_121_T_3[6:0] ? myVec_109 : _GEN_1046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1048 = 7'h6e == _myNewVec_121_T_3[6:0] ? myVec_110 : _GEN_1047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1049 = 7'h6f == _myNewVec_121_T_3[6:0] ? myVec_111 : _GEN_1048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1050 = 7'h70 == _myNewVec_121_T_3[6:0] ? myVec_112 : _GEN_1049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1051 = 7'h71 == _myNewVec_121_T_3[6:0] ? myVec_113 : _GEN_1050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1052 = 7'h72 == _myNewVec_121_T_3[6:0] ? myVec_114 : _GEN_1051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1053 = 7'h73 == _myNewVec_121_T_3[6:0] ? myVec_115 : _GEN_1052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1054 = 7'h74 == _myNewVec_121_T_3[6:0] ? myVec_116 : _GEN_1053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1055 = 7'h75 == _myNewVec_121_T_3[6:0] ? myVec_117 : _GEN_1054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1056 = 7'h76 == _myNewVec_121_T_3[6:0] ? myVec_118 : _GEN_1055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1057 = 7'h77 == _myNewVec_121_T_3[6:0] ? myVec_119 : _GEN_1056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1058 = 7'h78 == _myNewVec_121_T_3[6:0] ? myVec_120 : _GEN_1057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1059 = 7'h79 == _myNewVec_121_T_3[6:0] ? myVec_121 : _GEN_1058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1060 = 7'h7a == _myNewVec_121_T_3[6:0] ? myVec_122 : _GEN_1059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1061 = 7'h7b == _myNewVec_121_T_3[6:0] ? myVec_123 : _GEN_1060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1062 = 7'h7c == _myNewVec_121_T_3[6:0] ? myVec_124 : _GEN_1061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1063 = 7'h7d == _myNewVec_121_T_3[6:0] ? myVec_125 : _GEN_1062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1064 = 7'h7e == _myNewVec_121_T_3[6:0] ? myVec_126 : _GEN_1063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_121 = 7'h7f == _myNewVec_121_T_3[6:0] ? myVec_127 : _GEN_1064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_120_T_3 = _myNewVec_127_T_1 + 16'h7; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1067 = 7'h1 == _myNewVec_120_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1068 = 7'h2 == _myNewVec_120_T_3[6:0] ? myVec_2 : _GEN_1067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1069 = 7'h3 == _myNewVec_120_T_3[6:0] ? myVec_3 : _GEN_1068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1070 = 7'h4 == _myNewVec_120_T_3[6:0] ? myVec_4 : _GEN_1069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1071 = 7'h5 == _myNewVec_120_T_3[6:0] ? myVec_5 : _GEN_1070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1072 = 7'h6 == _myNewVec_120_T_3[6:0] ? myVec_6 : _GEN_1071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1073 = 7'h7 == _myNewVec_120_T_3[6:0] ? myVec_7 : _GEN_1072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1074 = 7'h8 == _myNewVec_120_T_3[6:0] ? myVec_8 : _GEN_1073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1075 = 7'h9 == _myNewVec_120_T_3[6:0] ? myVec_9 : _GEN_1074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1076 = 7'ha == _myNewVec_120_T_3[6:0] ? myVec_10 : _GEN_1075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1077 = 7'hb == _myNewVec_120_T_3[6:0] ? myVec_11 : _GEN_1076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1078 = 7'hc == _myNewVec_120_T_3[6:0] ? myVec_12 : _GEN_1077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1079 = 7'hd == _myNewVec_120_T_3[6:0] ? myVec_13 : _GEN_1078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1080 = 7'he == _myNewVec_120_T_3[6:0] ? myVec_14 : _GEN_1079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1081 = 7'hf == _myNewVec_120_T_3[6:0] ? myVec_15 : _GEN_1080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1082 = 7'h10 == _myNewVec_120_T_3[6:0] ? myVec_16 : _GEN_1081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1083 = 7'h11 == _myNewVec_120_T_3[6:0] ? myVec_17 : _GEN_1082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1084 = 7'h12 == _myNewVec_120_T_3[6:0] ? myVec_18 : _GEN_1083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1085 = 7'h13 == _myNewVec_120_T_3[6:0] ? myVec_19 : _GEN_1084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1086 = 7'h14 == _myNewVec_120_T_3[6:0] ? myVec_20 : _GEN_1085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1087 = 7'h15 == _myNewVec_120_T_3[6:0] ? myVec_21 : _GEN_1086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1088 = 7'h16 == _myNewVec_120_T_3[6:0] ? myVec_22 : _GEN_1087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1089 = 7'h17 == _myNewVec_120_T_3[6:0] ? myVec_23 : _GEN_1088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1090 = 7'h18 == _myNewVec_120_T_3[6:0] ? myVec_24 : _GEN_1089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1091 = 7'h19 == _myNewVec_120_T_3[6:0] ? myVec_25 : _GEN_1090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1092 = 7'h1a == _myNewVec_120_T_3[6:0] ? myVec_26 : _GEN_1091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1093 = 7'h1b == _myNewVec_120_T_3[6:0] ? myVec_27 : _GEN_1092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1094 = 7'h1c == _myNewVec_120_T_3[6:0] ? myVec_28 : _GEN_1093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1095 = 7'h1d == _myNewVec_120_T_3[6:0] ? myVec_29 : _GEN_1094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1096 = 7'h1e == _myNewVec_120_T_3[6:0] ? myVec_30 : _GEN_1095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1097 = 7'h1f == _myNewVec_120_T_3[6:0] ? myVec_31 : _GEN_1096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1098 = 7'h20 == _myNewVec_120_T_3[6:0] ? myVec_32 : _GEN_1097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1099 = 7'h21 == _myNewVec_120_T_3[6:0] ? myVec_33 : _GEN_1098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1100 = 7'h22 == _myNewVec_120_T_3[6:0] ? myVec_34 : _GEN_1099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1101 = 7'h23 == _myNewVec_120_T_3[6:0] ? myVec_35 : _GEN_1100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1102 = 7'h24 == _myNewVec_120_T_3[6:0] ? myVec_36 : _GEN_1101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1103 = 7'h25 == _myNewVec_120_T_3[6:0] ? myVec_37 : _GEN_1102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1104 = 7'h26 == _myNewVec_120_T_3[6:0] ? myVec_38 : _GEN_1103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1105 = 7'h27 == _myNewVec_120_T_3[6:0] ? myVec_39 : _GEN_1104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1106 = 7'h28 == _myNewVec_120_T_3[6:0] ? myVec_40 : _GEN_1105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1107 = 7'h29 == _myNewVec_120_T_3[6:0] ? myVec_41 : _GEN_1106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1108 = 7'h2a == _myNewVec_120_T_3[6:0] ? myVec_42 : _GEN_1107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1109 = 7'h2b == _myNewVec_120_T_3[6:0] ? myVec_43 : _GEN_1108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1110 = 7'h2c == _myNewVec_120_T_3[6:0] ? myVec_44 : _GEN_1109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1111 = 7'h2d == _myNewVec_120_T_3[6:0] ? myVec_45 : _GEN_1110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1112 = 7'h2e == _myNewVec_120_T_3[6:0] ? myVec_46 : _GEN_1111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1113 = 7'h2f == _myNewVec_120_T_3[6:0] ? myVec_47 : _GEN_1112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1114 = 7'h30 == _myNewVec_120_T_3[6:0] ? myVec_48 : _GEN_1113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1115 = 7'h31 == _myNewVec_120_T_3[6:0] ? myVec_49 : _GEN_1114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1116 = 7'h32 == _myNewVec_120_T_3[6:0] ? myVec_50 : _GEN_1115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1117 = 7'h33 == _myNewVec_120_T_3[6:0] ? myVec_51 : _GEN_1116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1118 = 7'h34 == _myNewVec_120_T_3[6:0] ? myVec_52 : _GEN_1117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1119 = 7'h35 == _myNewVec_120_T_3[6:0] ? myVec_53 : _GEN_1118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1120 = 7'h36 == _myNewVec_120_T_3[6:0] ? myVec_54 : _GEN_1119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1121 = 7'h37 == _myNewVec_120_T_3[6:0] ? myVec_55 : _GEN_1120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1122 = 7'h38 == _myNewVec_120_T_3[6:0] ? myVec_56 : _GEN_1121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1123 = 7'h39 == _myNewVec_120_T_3[6:0] ? myVec_57 : _GEN_1122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1124 = 7'h3a == _myNewVec_120_T_3[6:0] ? myVec_58 : _GEN_1123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1125 = 7'h3b == _myNewVec_120_T_3[6:0] ? myVec_59 : _GEN_1124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1126 = 7'h3c == _myNewVec_120_T_3[6:0] ? myVec_60 : _GEN_1125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1127 = 7'h3d == _myNewVec_120_T_3[6:0] ? myVec_61 : _GEN_1126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1128 = 7'h3e == _myNewVec_120_T_3[6:0] ? myVec_62 : _GEN_1127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1129 = 7'h3f == _myNewVec_120_T_3[6:0] ? myVec_63 : _GEN_1128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1130 = 7'h40 == _myNewVec_120_T_3[6:0] ? myVec_64 : _GEN_1129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1131 = 7'h41 == _myNewVec_120_T_3[6:0] ? myVec_65 : _GEN_1130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1132 = 7'h42 == _myNewVec_120_T_3[6:0] ? myVec_66 : _GEN_1131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1133 = 7'h43 == _myNewVec_120_T_3[6:0] ? myVec_67 : _GEN_1132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1134 = 7'h44 == _myNewVec_120_T_3[6:0] ? myVec_68 : _GEN_1133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1135 = 7'h45 == _myNewVec_120_T_3[6:0] ? myVec_69 : _GEN_1134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1136 = 7'h46 == _myNewVec_120_T_3[6:0] ? myVec_70 : _GEN_1135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1137 = 7'h47 == _myNewVec_120_T_3[6:0] ? myVec_71 : _GEN_1136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1138 = 7'h48 == _myNewVec_120_T_3[6:0] ? myVec_72 : _GEN_1137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1139 = 7'h49 == _myNewVec_120_T_3[6:0] ? myVec_73 : _GEN_1138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1140 = 7'h4a == _myNewVec_120_T_3[6:0] ? myVec_74 : _GEN_1139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1141 = 7'h4b == _myNewVec_120_T_3[6:0] ? myVec_75 : _GEN_1140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1142 = 7'h4c == _myNewVec_120_T_3[6:0] ? myVec_76 : _GEN_1141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1143 = 7'h4d == _myNewVec_120_T_3[6:0] ? myVec_77 : _GEN_1142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1144 = 7'h4e == _myNewVec_120_T_3[6:0] ? myVec_78 : _GEN_1143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1145 = 7'h4f == _myNewVec_120_T_3[6:0] ? myVec_79 : _GEN_1144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1146 = 7'h50 == _myNewVec_120_T_3[6:0] ? myVec_80 : _GEN_1145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1147 = 7'h51 == _myNewVec_120_T_3[6:0] ? myVec_81 : _GEN_1146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1148 = 7'h52 == _myNewVec_120_T_3[6:0] ? myVec_82 : _GEN_1147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1149 = 7'h53 == _myNewVec_120_T_3[6:0] ? myVec_83 : _GEN_1148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1150 = 7'h54 == _myNewVec_120_T_3[6:0] ? myVec_84 : _GEN_1149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1151 = 7'h55 == _myNewVec_120_T_3[6:0] ? myVec_85 : _GEN_1150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1152 = 7'h56 == _myNewVec_120_T_3[6:0] ? myVec_86 : _GEN_1151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1153 = 7'h57 == _myNewVec_120_T_3[6:0] ? myVec_87 : _GEN_1152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1154 = 7'h58 == _myNewVec_120_T_3[6:0] ? myVec_88 : _GEN_1153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1155 = 7'h59 == _myNewVec_120_T_3[6:0] ? myVec_89 : _GEN_1154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1156 = 7'h5a == _myNewVec_120_T_3[6:0] ? myVec_90 : _GEN_1155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1157 = 7'h5b == _myNewVec_120_T_3[6:0] ? myVec_91 : _GEN_1156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1158 = 7'h5c == _myNewVec_120_T_3[6:0] ? myVec_92 : _GEN_1157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1159 = 7'h5d == _myNewVec_120_T_3[6:0] ? myVec_93 : _GEN_1158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1160 = 7'h5e == _myNewVec_120_T_3[6:0] ? myVec_94 : _GEN_1159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1161 = 7'h5f == _myNewVec_120_T_3[6:0] ? myVec_95 : _GEN_1160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1162 = 7'h60 == _myNewVec_120_T_3[6:0] ? myVec_96 : _GEN_1161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1163 = 7'h61 == _myNewVec_120_T_3[6:0] ? myVec_97 : _GEN_1162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1164 = 7'h62 == _myNewVec_120_T_3[6:0] ? myVec_98 : _GEN_1163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1165 = 7'h63 == _myNewVec_120_T_3[6:0] ? myVec_99 : _GEN_1164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1166 = 7'h64 == _myNewVec_120_T_3[6:0] ? myVec_100 : _GEN_1165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1167 = 7'h65 == _myNewVec_120_T_3[6:0] ? myVec_101 : _GEN_1166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1168 = 7'h66 == _myNewVec_120_T_3[6:0] ? myVec_102 : _GEN_1167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1169 = 7'h67 == _myNewVec_120_T_3[6:0] ? myVec_103 : _GEN_1168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1170 = 7'h68 == _myNewVec_120_T_3[6:0] ? myVec_104 : _GEN_1169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1171 = 7'h69 == _myNewVec_120_T_3[6:0] ? myVec_105 : _GEN_1170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1172 = 7'h6a == _myNewVec_120_T_3[6:0] ? myVec_106 : _GEN_1171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1173 = 7'h6b == _myNewVec_120_T_3[6:0] ? myVec_107 : _GEN_1172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1174 = 7'h6c == _myNewVec_120_T_3[6:0] ? myVec_108 : _GEN_1173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1175 = 7'h6d == _myNewVec_120_T_3[6:0] ? myVec_109 : _GEN_1174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1176 = 7'h6e == _myNewVec_120_T_3[6:0] ? myVec_110 : _GEN_1175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1177 = 7'h6f == _myNewVec_120_T_3[6:0] ? myVec_111 : _GEN_1176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1178 = 7'h70 == _myNewVec_120_T_3[6:0] ? myVec_112 : _GEN_1177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1179 = 7'h71 == _myNewVec_120_T_3[6:0] ? myVec_113 : _GEN_1178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1180 = 7'h72 == _myNewVec_120_T_3[6:0] ? myVec_114 : _GEN_1179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1181 = 7'h73 == _myNewVec_120_T_3[6:0] ? myVec_115 : _GEN_1180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1182 = 7'h74 == _myNewVec_120_T_3[6:0] ? myVec_116 : _GEN_1181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1183 = 7'h75 == _myNewVec_120_T_3[6:0] ? myVec_117 : _GEN_1182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1184 = 7'h76 == _myNewVec_120_T_3[6:0] ? myVec_118 : _GEN_1183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1185 = 7'h77 == _myNewVec_120_T_3[6:0] ? myVec_119 : _GEN_1184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1186 = 7'h78 == _myNewVec_120_T_3[6:0] ? myVec_120 : _GEN_1185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1187 = 7'h79 == _myNewVec_120_T_3[6:0] ? myVec_121 : _GEN_1186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1188 = 7'h7a == _myNewVec_120_T_3[6:0] ? myVec_122 : _GEN_1187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1189 = 7'h7b == _myNewVec_120_T_3[6:0] ? myVec_123 : _GEN_1188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1190 = 7'h7c == _myNewVec_120_T_3[6:0] ? myVec_124 : _GEN_1189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1191 = 7'h7d == _myNewVec_120_T_3[6:0] ? myVec_125 : _GEN_1190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1192 = 7'h7e == _myNewVec_120_T_3[6:0] ? myVec_126 : _GEN_1191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_120 = 7'h7f == _myNewVec_120_T_3[6:0] ? myVec_127 : _GEN_1192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_119_T_3 = _myNewVec_127_T_1 + 16'h8; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1195 = 7'h1 == _myNewVec_119_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1196 = 7'h2 == _myNewVec_119_T_3[6:0] ? myVec_2 : _GEN_1195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1197 = 7'h3 == _myNewVec_119_T_3[6:0] ? myVec_3 : _GEN_1196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1198 = 7'h4 == _myNewVec_119_T_3[6:0] ? myVec_4 : _GEN_1197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1199 = 7'h5 == _myNewVec_119_T_3[6:0] ? myVec_5 : _GEN_1198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1200 = 7'h6 == _myNewVec_119_T_3[6:0] ? myVec_6 : _GEN_1199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1201 = 7'h7 == _myNewVec_119_T_3[6:0] ? myVec_7 : _GEN_1200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1202 = 7'h8 == _myNewVec_119_T_3[6:0] ? myVec_8 : _GEN_1201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1203 = 7'h9 == _myNewVec_119_T_3[6:0] ? myVec_9 : _GEN_1202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1204 = 7'ha == _myNewVec_119_T_3[6:0] ? myVec_10 : _GEN_1203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1205 = 7'hb == _myNewVec_119_T_3[6:0] ? myVec_11 : _GEN_1204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1206 = 7'hc == _myNewVec_119_T_3[6:0] ? myVec_12 : _GEN_1205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1207 = 7'hd == _myNewVec_119_T_3[6:0] ? myVec_13 : _GEN_1206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1208 = 7'he == _myNewVec_119_T_3[6:0] ? myVec_14 : _GEN_1207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1209 = 7'hf == _myNewVec_119_T_3[6:0] ? myVec_15 : _GEN_1208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1210 = 7'h10 == _myNewVec_119_T_3[6:0] ? myVec_16 : _GEN_1209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1211 = 7'h11 == _myNewVec_119_T_3[6:0] ? myVec_17 : _GEN_1210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1212 = 7'h12 == _myNewVec_119_T_3[6:0] ? myVec_18 : _GEN_1211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1213 = 7'h13 == _myNewVec_119_T_3[6:0] ? myVec_19 : _GEN_1212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1214 = 7'h14 == _myNewVec_119_T_3[6:0] ? myVec_20 : _GEN_1213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1215 = 7'h15 == _myNewVec_119_T_3[6:0] ? myVec_21 : _GEN_1214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1216 = 7'h16 == _myNewVec_119_T_3[6:0] ? myVec_22 : _GEN_1215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1217 = 7'h17 == _myNewVec_119_T_3[6:0] ? myVec_23 : _GEN_1216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1218 = 7'h18 == _myNewVec_119_T_3[6:0] ? myVec_24 : _GEN_1217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1219 = 7'h19 == _myNewVec_119_T_3[6:0] ? myVec_25 : _GEN_1218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1220 = 7'h1a == _myNewVec_119_T_3[6:0] ? myVec_26 : _GEN_1219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1221 = 7'h1b == _myNewVec_119_T_3[6:0] ? myVec_27 : _GEN_1220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1222 = 7'h1c == _myNewVec_119_T_3[6:0] ? myVec_28 : _GEN_1221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1223 = 7'h1d == _myNewVec_119_T_3[6:0] ? myVec_29 : _GEN_1222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1224 = 7'h1e == _myNewVec_119_T_3[6:0] ? myVec_30 : _GEN_1223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1225 = 7'h1f == _myNewVec_119_T_3[6:0] ? myVec_31 : _GEN_1224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1226 = 7'h20 == _myNewVec_119_T_3[6:0] ? myVec_32 : _GEN_1225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1227 = 7'h21 == _myNewVec_119_T_3[6:0] ? myVec_33 : _GEN_1226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1228 = 7'h22 == _myNewVec_119_T_3[6:0] ? myVec_34 : _GEN_1227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1229 = 7'h23 == _myNewVec_119_T_3[6:0] ? myVec_35 : _GEN_1228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1230 = 7'h24 == _myNewVec_119_T_3[6:0] ? myVec_36 : _GEN_1229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1231 = 7'h25 == _myNewVec_119_T_3[6:0] ? myVec_37 : _GEN_1230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1232 = 7'h26 == _myNewVec_119_T_3[6:0] ? myVec_38 : _GEN_1231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1233 = 7'h27 == _myNewVec_119_T_3[6:0] ? myVec_39 : _GEN_1232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1234 = 7'h28 == _myNewVec_119_T_3[6:0] ? myVec_40 : _GEN_1233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1235 = 7'h29 == _myNewVec_119_T_3[6:0] ? myVec_41 : _GEN_1234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1236 = 7'h2a == _myNewVec_119_T_3[6:0] ? myVec_42 : _GEN_1235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1237 = 7'h2b == _myNewVec_119_T_3[6:0] ? myVec_43 : _GEN_1236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1238 = 7'h2c == _myNewVec_119_T_3[6:0] ? myVec_44 : _GEN_1237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1239 = 7'h2d == _myNewVec_119_T_3[6:0] ? myVec_45 : _GEN_1238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1240 = 7'h2e == _myNewVec_119_T_3[6:0] ? myVec_46 : _GEN_1239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1241 = 7'h2f == _myNewVec_119_T_3[6:0] ? myVec_47 : _GEN_1240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1242 = 7'h30 == _myNewVec_119_T_3[6:0] ? myVec_48 : _GEN_1241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1243 = 7'h31 == _myNewVec_119_T_3[6:0] ? myVec_49 : _GEN_1242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1244 = 7'h32 == _myNewVec_119_T_3[6:0] ? myVec_50 : _GEN_1243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1245 = 7'h33 == _myNewVec_119_T_3[6:0] ? myVec_51 : _GEN_1244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1246 = 7'h34 == _myNewVec_119_T_3[6:0] ? myVec_52 : _GEN_1245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1247 = 7'h35 == _myNewVec_119_T_3[6:0] ? myVec_53 : _GEN_1246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1248 = 7'h36 == _myNewVec_119_T_3[6:0] ? myVec_54 : _GEN_1247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1249 = 7'h37 == _myNewVec_119_T_3[6:0] ? myVec_55 : _GEN_1248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1250 = 7'h38 == _myNewVec_119_T_3[6:0] ? myVec_56 : _GEN_1249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1251 = 7'h39 == _myNewVec_119_T_3[6:0] ? myVec_57 : _GEN_1250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1252 = 7'h3a == _myNewVec_119_T_3[6:0] ? myVec_58 : _GEN_1251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1253 = 7'h3b == _myNewVec_119_T_3[6:0] ? myVec_59 : _GEN_1252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1254 = 7'h3c == _myNewVec_119_T_3[6:0] ? myVec_60 : _GEN_1253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1255 = 7'h3d == _myNewVec_119_T_3[6:0] ? myVec_61 : _GEN_1254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1256 = 7'h3e == _myNewVec_119_T_3[6:0] ? myVec_62 : _GEN_1255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1257 = 7'h3f == _myNewVec_119_T_3[6:0] ? myVec_63 : _GEN_1256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1258 = 7'h40 == _myNewVec_119_T_3[6:0] ? myVec_64 : _GEN_1257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1259 = 7'h41 == _myNewVec_119_T_3[6:0] ? myVec_65 : _GEN_1258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1260 = 7'h42 == _myNewVec_119_T_3[6:0] ? myVec_66 : _GEN_1259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1261 = 7'h43 == _myNewVec_119_T_3[6:0] ? myVec_67 : _GEN_1260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1262 = 7'h44 == _myNewVec_119_T_3[6:0] ? myVec_68 : _GEN_1261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1263 = 7'h45 == _myNewVec_119_T_3[6:0] ? myVec_69 : _GEN_1262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1264 = 7'h46 == _myNewVec_119_T_3[6:0] ? myVec_70 : _GEN_1263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1265 = 7'h47 == _myNewVec_119_T_3[6:0] ? myVec_71 : _GEN_1264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1266 = 7'h48 == _myNewVec_119_T_3[6:0] ? myVec_72 : _GEN_1265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1267 = 7'h49 == _myNewVec_119_T_3[6:0] ? myVec_73 : _GEN_1266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1268 = 7'h4a == _myNewVec_119_T_3[6:0] ? myVec_74 : _GEN_1267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1269 = 7'h4b == _myNewVec_119_T_3[6:0] ? myVec_75 : _GEN_1268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1270 = 7'h4c == _myNewVec_119_T_3[6:0] ? myVec_76 : _GEN_1269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1271 = 7'h4d == _myNewVec_119_T_3[6:0] ? myVec_77 : _GEN_1270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1272 = 7'h4e == _myNewVec_119_T_3[6:0] ? myVec_78 : _GEN_1271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1273 = 7'h4f == _myNewVec_119_T_3[6:0] ? myVec_79 : _GEN_1272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1274 = 7'h50 == _myNewVec_119_T_3[6:0] ? myVec_80 : _GEN_1273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1275 = 7'h51 == _myNewVec_119_T_3[6:0] ? myVec_81 : _GEN_1274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1276 = 7'h52 == _myNewVec_119_T_3[6:0] ? myVec_82 : _GEN_1275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1277 = 7'h53 == _myNewVec_119_T_3[6:0] ? myVec_83 : _GEN_1276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1278 = 7'h54 == _myNewVec_119_T_3[6:0] ? myVec_84 : _GEN_1277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1279 = 7'h55 == _myNewVec_119_T_3[6:0] ? myVec_85 : _GEN_1278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1280 = 7'h56 == _myNewVec_119_T_3[6:0] ? myVec_86 : _GEN_1279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1281 = 7'h57 == _myNewVec_119_T_3[6:0] ? myVec_87 : _GEN_1280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1282 = 7'h58 == _myNewVec_119_T_3[6:0] ? myVec_88 : _GEN_1281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1283 = 7'h59 == _myNewVec_119_T_3[6:0] ? myVec_89 : _GEN_1282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1284 = 7'h5a == _myNewVec_119_T_3[6:0] ? myVec_90 : _GEN_1283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1285 = 7'h5b == _myNewVec_119_T_3[6:0] ? myVec_91 : _GEN_1284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1286 = 7'h5c == _myNewVec_119_T_3[6:0] ? myVec_92 : _GEN_1285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1287 = 7'h5d == _myNewVec_119_T_3[6:0] ? myVec_93 : _GEN_1286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1288 = 7'h5e == _myNewVec_119_T_3[6:0] ? myVec_94 : _GEN_1287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1289 = 7'h5f == _myNewVec_119_T_3[6:0] ? myVec_95 : _GEN_1288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1290 = 7'h60 == _myNewVec_119_T_3[6:0] ? myVec_96 : _GEN_1289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1291 = 7'h61 == _myNewVec_119_T_3[6:0] ? myVec_97 : _GEN_1290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1292 = 7'h62 == _myNewVec_119_T_3[6:0] ? myVec_98 : _GEN_1291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1293 = 7'h63 == _myNewVec_119_T_3[6:0] ? myVec_99 : _GEN_1292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1294 = 7'h64 == _myNewVec_119_T_3[6:0] ? myVec_100 : _GEN_1293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1295 = 7'h65 == _myNewVec_119_T_3[6:0] ? myVec_101 : _GEN_1294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1296 = 7'h66 == _myNewVec_119_T_3[6:0] ? myVec_102 : _GEN_1295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1297 = 7'h67 == _myNewVec_119_T_3[6:0] ? myVec_103 : _GEN_1296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1298 = 7'h68 == _myNewVec_119_T_3[6:0] ? myVec_104 : _GEN_1297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1299 = 7'h69 == _myNewVec_119_T_3[6:0] ? myVec_105 : _GEN_1298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1300 = 7'h6a == _myNewVec_119_T_3[6:0] ? myVec_106 : _GEN_1299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1301 = 7'h6b == _myNewVec_119_T_3[6:0] ? myVec_107 : _GEN_1300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1302 = 7'h6c == _myNewVec_119_T_3[6:0] ? myVec_108 : _GEN_1301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1303 = 7'h6d == _myNewVec_119_T_3[6:0] ? myVec_109 : _GEN_1302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1304 = 7'h6e == _myNewVec_119_T_3[6:0] ? myVec_110 : _GEN_1303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1305 = 7'h6f == _myNewVec_119_T_3[6:0] ? myVec_111 : _GEN_1304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1306 = 7'h70 == _myNewVec_119_T_3[6:0] ? myVec_112 : _GEN_1305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1307 = 7'h71 == _myNewVec_119_T_3[6:0] ? myVec_113 : _GEN_1306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1308 = 7'h72 == _myNewVec_119_T_3[6:0] ? myVec_114 : _GEN_1307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1309 = 7'h73 == _myNewVec_119_T_3[6:0] ? myVec_115 : _GEN_1308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1310 = 7'h74 == _myNewVec_119_T_3[6:0] ? myVec_116 : _GEN_1309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1311 = 7'h75 == _myNewVec_119_T_3[6:0] ? myVec_117 : _GEN_1310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1312 = 7'h76 == _myNewVec_119_T_3[6:0] ? myVec_118 : _GEN_1311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1313 = 7'h77 == _myNewVec_119_T_3[6:0] ? myVec_119 : _GEN_1312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1314 = 7'h78 == _myNewVec_119_T_3[6:0] ? myVec_120 : _GEN_1313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1315 = 7'h79 == _myNewVec_119_T_3[6:0] ? myVec_121 : _GEN_1314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1316 = 7'h7a == _myNewVec_119_T_3[6:0] ? myVec_122 : _GEN_1315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1317 = 7'h7b == _myNewVec_119_T_3[6:0] ? myVec_123 : _GEN_1316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1318 = 7'h7c == _myNewVec_119_T_3[6:0] ? myVec_124 : _GEN_1317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1319 = 7'h7d == _myNewVec_119_T_3[6:0] ? myVec_125 : _GEN_1318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1320 = 7'h7e == _myNewVec_119_T_3[6:0] ? myVec_126 : _GEN_1319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_119 = 7'h7f == _myNewVec_119_T_3[6:0] ? myVec_127 : _GEN_1320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_118_T_3 = _myNewVec_127_T_1 + 16'h9; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1323 = 7'h1 == _myNewVec_118_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1324 = 7'h2 == _myNewVec_118_T_3[6:0] ? myVec_2 : _GEN_1323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1325 = 7'h3 == _myNewVec_118_T_3[6:0] ? myVec_3 : _GEN_1324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1326 = 7'h4 == _myNewVec_118_T_3[6:0] ? myVec_4 : _GEN_1325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1327 = 7'h5 == _myNewVec_118_T_3[6:0] ? myVec_5 : _GEN_1326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1328 = 7'h6 == _myNewVec_118_T_3[6:0] ? myVec_6 : _GEN_1327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1329 = 7'h7 == _myNewVec_118_T_3[6:0] ? myVec_7 : _GEN_1328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1330 = 7'h8 == _myNewVec_118_T_3[6:0] ? myVec_8 : _GEN_1329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1331 = 7'h9 == _myNewVec_118_T_3[6:0] ? myVec_9 : _GEN_1330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1332 = 7'ha == _myNewVec_118_T_3[6:0] ? myVec_10 : _GEN_1331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1333 = 7'hb == _myNewVec_118_T_3[6:0] ? myVec_11 : _GEN_1332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1334 = 7'hc == _myNewVec_118_T_3[6:0] ? myVec_12 : _GEN_1333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1335 = 7'hd == _myNewVec_118_T_3[6:0] ? myVec_13 : _GEN_1334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1336 = 7'he == _myNewVec_118_T_3[6:0] ? myVec_14 : _GEN_1335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1337 = 7'hf == _myNewVec_118_T_3[6:0] ? myVec_15 : _GEN_1336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1338 = 7'h10 == _myNewVec_118_T_3[6:0] ? myVec_16 : _GEN_1337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1339 = 7'h11 == _myNewVec_118_T_3[6:0] ? myVec_17 : _GEN_1338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1340 = 7'h12 == _myNewVec_118_T_3[6:0] ? myVec_18 : _GEN_1339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1341 = 7'h13 == _myNewVec_118_T_3[6:0] ? myVec_19 : _GEN_1340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1342 = 7'h14 == _myNewVec_118_T_3[6:0] ? myVec_20 : _GEN_1341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1343 = 7'h15 == _myNewVec_118_T_3[6:0] ? myVec_21 : _GEN_1342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1344 = 7'h16 == _myNewVec_118_T_3[6:0] ? myVec_22 : _GEN_1343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1345 = 7'h17 == _myNewVec_118_T_3[6:0] ? myVec_23 : _GEN_1344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1346 = 7'h18 == _myNewVec_118_T_3[6:0] ? myVec_24 : _GEN_1345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1347 = 7'h19 == _myNewVec_118_T_3[6:0] ? myVec_25 : _GEN_1346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1348 = 7'h1a == _myNewVec_118_T_3[6:0] ? myVec_26 : _GEN_1347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1349 = 7'h1b == _myNewVec_118_T_3[6:0] ? myVec_27 : _GEN_1348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1350 = 7'h1c == _myNewVec_118_T_3[6:0] ? myVec_28 : _GEN_1349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1351 = 7'h1d == _myNewVec_118_T_3[6:0] ? myVec_29 : _GEN_1350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1352 = 7'h1e == _myNewVec_118_T_3[6:0] ? myVec_30 : _GEN_1351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1353 = 7'h1f == _myNewVec_118_T_3[6:0] ? myVec_31 : _GEN_1352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1354 = 7'h20 == _myNewVec_118_T_3[6:0] ? myVec_32 : _GEN_1353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1355 = 7'h21 == _myNewVec_118_T_3[6:0] ? myVec_33 : _GEN_1354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1356 = 7'h22 == _myNewVec_118_T_3[6:0] ? myVec_34 : _GEN_1355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1357 = 7'h23 == _myNewVec_118_T_3[6:0] ? myVec_35 : _GEN_1356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1358 = 7'h24 == _myNewVec_118_T_3[6:0] ? myVec_36 : _GEN_1357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1359 = 7'h25 == _myNewVec_118_T_3[6:0] ? myVec_37 : _GEN_1358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1360 = 7'h26 == _myNewVec_118_T_3[6:0] ? myVec_38 : _GEN_1359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1361 = 7'h27 == _myNewVec_118_T_3[6:0] ? myVec_39 : _GEN_1360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1362 = 7'h28 == _myNewVec_118_T_3[6:0] ? myVec_40 : _GEN_1361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1363 = 7'h29 == _myNewVec_118_T_3[6:0] ? myVec_41 : _GEN_1362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1364 = 7'h2a == _myNewVec_118_T_3[6:0] ? myVec_42 : _GEN_1363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1365 = 7'h2b == _myNewVec_118_T_3[6:0] ? myVec_43 : _GEN_1364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1366 = 7'h2c == _myNewVec_118_T_3[6:0] ? myVec_44 : _GEN_1365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1367 = 7'h2d == _myNewVec_118_T_3[6:0] ? myVec_45 : _GEN_1366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1368 = 7'h2e == _myNewVec_118_T_3[6:0] ? myVec_46 : _GEN_1367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1369 = 7'h2f == _myNewVec_118_T_3[6:0] ? myVec_47 : _GEN_1368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1370 = 7'h30 == _myNewVec_118_T_3[6:0] ? myVec_48 : _GEN_1369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1371 = 7'h31 == _myNewVec_118_T_3[6:0] ? myVec_49 : _GEN_1370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1372 = 7'h32 == _myNewVec_118_T_3[6:0] ? myVec_50 : _GEN_1371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1373 = 7'h33 == _myNewVec_118_T_3[6:0] ? myVec_51 : _GEN_1372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1374 = 7'h34 == _myNewVec_118_T_3[6:0] ? myVec_52 : _GEN_1373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1375 = 7'h35 == _myNewVec_118_T_3[6:0] ? myVec_53 : _GEN_1374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1376 = 7'h36 == _myNewVec_118_T_3[6:0] ? myVec_54 : _GEN_1375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1377 = 7'h37 == _myNewVec_118_T_3[6:0] ? myVec_55 : _GEN_1376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1378 = 7'h38 == _myNewVec_118_T_3[6:0] ? myVec_56 : _GEN_1377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1379 = 7'h39 == _myNewVec_118_T_3[6:0] ? myVec_57 : _GEN_1378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1380 = 7'h3a == _myNewVec_118_T_3[6:0] ? myVec_58 : _GEN_1379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1381 = 7'h3b == _myNewVec_118_T_3[6:0] ? myVec_59 : _GEN_1380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1382 = 7'h3c == _myNewVec_118_T_3[6:0] ? myVec_60 : _GEN_1381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1383 = 7'h3d == _myNewVec_118_T_3[6:0] ? myVec_61 : _GEN_1382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1384 = 7'h3e == _myNewVec_118_T_3[6:0] ? myVec_62 : _GEN_1383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1385 = 7'h3f == _myNewVec_118_T_3[6:0] ? myVec_63 : _GEN_1384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1386 = 7'h40 == _myNewVec_118_T_3[6:0] ? myVec_64 : _GEN_1385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1387 = 7'h41 == _myNewVec_118_T_3[6:0] ? myVec_65 : _GEN_1386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1388 = 7'h42 == _myNewVec_118_T_3[6:0] ? myVec_66 : _GEN_1387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1389 = 7'h43 == _myNewVec_118_T_3[6:0] ? myVec_67 : _GEN_1388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1390 = 7'h44 == _myNewVec_118_T_3[6:0] ? myVec_68 : _GEN_1389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1391 = 7'h45 == _myNewVec_118_T_3[6:0] ? myVec_69 : _GEN_1390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1392 = 7'h46 == _myNewVec_118_T_3[6:0] ? myVec_70 : _GEN_1391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1393 = 7'h47 == _myNewVec_118_T_3[6:0] ? myVec_71 : _GEN_1392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1394 = 7'h48 == _myNewVec_118_T_3[6:0] ? myVec_72 : _GEN_1393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1395 = 7'h49 == _myNewVec_118_T_3[6:0] ? myVec_73 : _GEN_1394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1396 = 7'h4a == _myNewVec_118_T_3[6:0] ? myVec_74 : _GEN_1395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1397 = 7'h4b == _myNewVec_118_T_3[6:0] ? myVec_75 : _GEN_1396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1398 = 7'h4c == _myNewVec_118_T_3[6:0] ? myVec_76 : _GEN_1397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1399 = 7'h4d == _myNewVec_118_T_3[6:0] ? myVec_77 : _GEN_1398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1400 = 7'h4e == _myNewVec_118_T_3[6:0] ? myVec_78 : _GEN_1399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1401 = 7'h4f == _myNewVec_118_T_3[6:0] ? myVec_79 : _GEN_1400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1402 = 7'h50 == _myNewVec_118_T_3[6:0] ? myVec_80 : _GEN_1401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1403 = 7'h51 == _myNewVec_118_T_3[6:0] ? myVec_81 : _GEN_1402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1404 = 7'h52 == _myNewVec_118_T_3[6:0] ? myVec_82 : _GEN_1403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1405 = 7'h53 == _myNewVec_118_T_3[6:0] ? myVec_83 : _GEN_1404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1406 = 7'h54 == _myNewVec_118_T_3[6:0] ? myVec_84 : _GEN_1405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1407 = 7'h55 == _myNewVec_118_T_3[6:0] ? myVec_85 : _GEN_1406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1408 = 7'h56 == _myNewVec_118_T_3[6:0] ? myVec_86 : _GEN_1407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1409 = 7'h57 == _myNewVec_118_T_3[6:0] ? myVec_87 : _GEN_1408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1410 = 7'h58 == _myNewVec_118_T_3[6:0] ? myVec_88 : _GEN_1409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1411 = 7'h59 == _myNewVec_118_T_3[6:0] ? myVec_89 : _GEN_1410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1412 = 7'h5a == _myNewVec_118_T_3[6:0] ? myVec_90 : _GEN_1411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1413 = 7'h5b == _myNewVec_118_T_3[6:0] ? myVec_91 : _GEN_1412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1414 = 7'h5c == _myNewVec_118_T_3[6:0] ? myVec_92 : _GEN_1413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1415 = 7'h5d == _myNewVec_118_T_3[6:0] ? myVec_93 : _GEN_1414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1416 = 7'h5e == _myNewVec_118_T_3[6:0] ? myVec_94 : _GEN_1415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1417 = 7'h5f == _myNewVec_118_T_3[6:0] ? myVec_95 : _GEN_1416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1418 = 7'h60 == _myNewVec_118_T_3[6:0] ? myVec_96 : _GEN_1417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1419 = 7'h61 == _myNewVec_118_T_3[6:0] ? myVec_97 : _GEN_1418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1420 = 7'h62 == _myNewVec_118_T_3[6:0] ? myVec_98 : _GEN_1419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1421 = 7'h63 == _myNewVec_118_T_3[6:0] ? myVec_99 : _GEN_1420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1422 = 7'h64 == _myNewVec_118_T_3[6:0] ? myVec_100 : _GEN_1421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1423 = 7'h65 == _myNewVec_118_T_3[6:0] ? myVec_101 : _GEN_1422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1424 = 7'h66 == _myNewVec_118_T_3[6:0] ? myVec_102 : _GEN_1423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1425 = 7'h67 == _myNewVec_118_T_3[6:0] ? myVec_103 : _GEN_1424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1426 = 7'h68 == _myNewVec_118_T_3[6:0] ? myVec_104 : _GEN_1425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1427 = 7'h69 == _myNewVec_118_T_3[6:0] ? myVec_105 : _GEN_1426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1428 = 7'h6a == _myNewVec_118_T_3[6:0] ? myVec_106 : _GEN_1427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1429 = 7'h6b == _myNewVec_118_T_3[6:0] ? myVec_107 : _GEN_1428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1430 = 7'h6c == _myNewVec_118_T_3[6:0] ? myVec_108 : _GEN_1429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1431 = 7'h6d == _myNewVec_118_T_3[6:0] ? myVec_109 : _GEN_1430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1432 = 7'h6e == _myNewVec_118_T_3[6:0] ? myVec_110 : _GEN_1431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1433 = 7'h6f == _myNewVec_118_T_3[6:0] ? myVec_111 : _GEN_1432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1434 = 7'h70 == _myNewVec_118_T_3[6:0] ? myVec_112 : _GEN_1433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1435 = 7'h71 == _myNewVec_118_T_3[6:0] ? myVec_113 : _GEN_1434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1436 = 7'h72 == _myNewVec_118_T_3[6:0] ? myVec_114 : _GEN_1435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1437 = 7'h73 == _myNewVec_118_T_3[6:0] ? myVec_115 : _GEN_1436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1438 = 7'h74 == _myNewVec_118_T_3[6:0] ? myVec_116 : _GEN_1437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1439 = 7'h75 == _myNewVec_118_T_3[6:0] ? myVec_117 : _GEN_1438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1440 = 7'h76 == _myNewVec_118_T_3[6:0] ? myVec_118 : _GEN_1439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1441 = 7'h77 == _myNewVec_118_T_3[6:0] ? myVec_119 : _GEN_1440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1442 = 7'h78 == _myNewVec_118_T_3[6:0] ? myVec_120 : _GEN_1441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1443 = 7'h79 == _myNewVec_118_T_3[6:0] ? myVec_121 : _GEN_1442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1444 = 7'h7a == _myNewVec_118_T_3[6:0] ? myVec_122 : _GEN_1443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1445 = 7'h7b == _myNewVec_118_T_3[6:0] ? myVec_123 : _GEN_1444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1446 = 7'h7c == _myNewVec_118_T_3[6:0] ? myVec_124 : _GEN_1445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1447 = 7'h7d == _myNewVec_118_T_3[6:0] ? myVec_125 : _GEN_1446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1448 = 7'h7e == _myNewVec_118_T_3[6:0] ? myVec_126 : _GEN_1447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_118 = 7'h7f == _myNewVec_118_T_3[6:0] ? myVec_127 : _GEN_1448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_117_T_3 = _myNewVec_127_T_1 + 16'ha; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1451 = 7'h1 == _myNewVec_117_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1452 = 7'h2 == _myNewVec_117_T_3[6:0] ? myVec_2 : _GEN_1451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1453 = 7'h3 == _myNewVec_117_T_3[6:0] ? myVec_3 : _GEN_1452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1454 = 7'h4 == _myNewVec_117_T_3[6:0] ? myVec_4 : _GEN_1453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1455 = 7'h5 == _myNewVec_117_T_3[6:0] ? myVec_5 : _GEN_1454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1456 = 7'h6 == _myNewVec_117_T_3[6:0] ? myVec_6 : _GEN_1455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1457 = 7'h7 == _myNewVec_117_T_3[6:0] ? myVec_7 : _GEN_1456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1458 = 7'h8 == _myNewVec_117_T_3[6:0] ? myVec_8 : _GEN_1457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1459 = 7'h9 == _myNewVec_117_T_3[6:0] ? myVec_9 : _GEN_1458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1460 = 7'ha == _myNewVec_117_T_3[6:0] ? myVec_10 : _GEN_1459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1461 = 7'hb == _myNewVec_117_T_3[6:0] ? myVec_11 : _GEN_1460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1462 = 7'hc == _myNewVec_117_T_3[6:0] ? myVec_12 : _GEN_1461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1463 = 7'hd == _myNewVec_117_T_3[6:0] ? myVec_13 : _GEN_1462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1464 = 7'he == _myNewVec_117_T_3[6:0] ? myVec_14 : _GEN_1463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1465 = 7'hf == _myNewVec_117_T_3[6:0] ? myVec_15 : _GEN_1464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1466 = 7'h10 == _myNewVec_117_T_3[6:0] ? myVec_16 : _GEN_1465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1467 = 7'h11 == _myNewVec_117_T_3[6:0] ? myVec_17 : _GEN_1466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1468 = 7'h12 == _myNewVec_117_T_3[6:0] ? myVec_18 : _GEN_1467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1469 = 7'h13 == _myNewVec_117_T_3[6:0] ? myVec_19 : _GEN_1468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1470 = 7'h14 == _myNewVec_117_T_3[6:0] ? myVec_20 : _GEN_1469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1471 = 7'h15 == _myNewVec_117_T_3[6:0] ? myVec_21 : _GEN_1470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1472 = 7'h16 == _myNewVec_117_T_3[6:0] ? myVec_22 : _GEN_1471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1473 = 7'h17 == _myNewVec_117_T_3[6:0] ? myVec_23 : _GEN_1472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1474 = 7'h18 == _myNewVec_117_T_3[6:0] ? myVec_24 : _GEN_1473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1475 = 7'h19 == _myNewVec_117_T_3[6:0] ? myVec_25 : _GEN_1474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1476 = 7'h1a == _myNewVec_117_T_3[6:0] ? myVec_26 : _GEN_1475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1477 = 7'h1b == _myNewVec_117_T_3[6:0] ? myVec_27 : _GEN_1476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1478 = 7'h1c == _myNewVec_117_T_3[6:0] ? myVec_28 : _GEN_1477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1479 = 7'h1d == _myNewVec_117_T_3[6:0] ? myVec_29 : _GEN_1478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1480 = 7'h1e == _myNewVec_117_T_3[6:0] ? myVec_30 : _GEN_1479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1481 = 7'h1f == _myNewVec_117_T_3[6:0] ? myVec_31 : _GEN_1480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1482 = 7'h20 == _myNewVec_117_T_3[6:0] ? myVec_32 : _GEN_1481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1483 = 7'h21 == _myNewVec_117_T_3[6:0] ? myVec_33 : _GEN_1482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1484 = 7'h22 == _myNewVec_117_T_3[6:0] ? myVec_34 : _GEN_1483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1485 = 7'h23 == _myNewVec_117_T_3[6:0] ? myVec_35 : _GEN_1484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1486 = 7'h24 == _myNewVec_117_T_3[6:0] ? myVec_36 : _GEN_1485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1487 = 7'h25 == _myNewVec_117_T_3[6:0] ? myVec_37 : _GEN_1486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1488 = 7'h26 == _myNewVec_117_T_3[6:0] ? myVec_38 : _GEN_1487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1489 = 7'h27 == _myNewVec_117_T_3[6:0] ? myVec_39 : _GEN_1488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1490 = 7'h28 == _myNewVec_117_T_3[6:0] ? myVec_40 : _GEN_1489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1491 = 7'h29 == _myNewVec_117_T_3[6:0] ? myVec_41 : _GEN_1490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1492 = 7'h2a == _myNewVec_117_T_3[6:0] ? myVec_42 : _GEN_1491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1493 = 7'h2b == _myNewVec_117_T_3[6:0] ? myVec_43 : _GEN_1492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1494 = 7'h2c == _myNewVec_117_T_3[6:0] ? myVec_44 : _GEN_1493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1495 = 7'h2d == _myNewVec_117_T_3[6:0] ? myVec_45 : _GEN_1494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1496 = 7'h2e == _myNewVec_117_T_3[6:0] ? myVec_46 : _GEN_1495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1497 = 7'h2f == _myNewVec_117_T_3[6:0] ? myVec_47 : _GEN_1496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1498 = 7'h30 == _myNewVec_117_T_3[6:0] ? myVec_48 : _GEN_1497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1499 = 7'h31 == _myNewVec_117_T_3[6:0] ? myVec_49 : _GEN_1498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1500 = 7'h32 == _myNewVec_117_T_3[6:0] ? myVec_50 : _GEN_1499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1501 = 7'h33 == _myNewVec_117_T_3[6:0] ? myVec_51 : _GEN_1500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1502 = 7'h34 == _myNewVec_117_T_3[6:0] ? myVec_52 : _GEN_1501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1503 = 7'h35 == _myNewVec_117_T_3[6:0] ? myVec_53 : _GEN_1502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1504 = 7'h36 == _myNewVec_117_T_3[6:0] ? myVec_54 : _GEN_1503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1505 = 7'h37 == _myNewVec_117_T_3[6:0] ? myVec_55 : _GEN_1504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1506 = 7'h38 == _myNewVec_117_T_3[6:0] ? myVec_56 : _GEN_1505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1507 = 7'h39 == _myNewVec_117_T_3[6:0] ? myVec_57 : _GEN_1506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1508 = 7'h3a == _myNewVec_117_T_3[6:0] ? myVec_58 : _GEN_1507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1509 = 7'h3b == _myNewVec_117_T_3[6:0] ? myVec_59 : _GEN_1508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1510 = 7'h3c == _myNewVec_117_T_3[6:0] ? myVec_60 : _GEN_1509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1511 = 7'h3d == _myNewVec_117_T_3[6:0] ? myVec_61 : _GEN_1510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1512 = 7'h3e == _myNewVec_117_T_3[6:0] ? myVec_62 : _GEN_1511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1513 = 7'h3f == _myNewVec_117_T_3[6:0] ? myVec_63 : _GEN_1512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1514 = 7'h40 == _myNewVec_117_T_3[6:0] ? myVec_64 : _GEN_1513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1515 = 7'h41 == _myNewVec_117_T_3[6:0] ? myVec_65 : _GEN_1514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1516 = 7'h42 == _myNewVec_117_T_3[6:0] ? myVec_66 : _GEN_1515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1517 = 7'h43 == _myNewVec_117_T_3[6:0] ? myVec_67 : _GEN_1516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1518 = 7'h44 == _myNewVec_117_T_3[6:0] ? myVec_68 : _GEN_1517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1519 = 7'h45 == _myNewVec_117_T_3[6:0] ? myVec_69 : _GEN_1518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1520 = 7'h46 == _myNewVec_117_T_3[6:0] ? myVec_70 : _GEN_1519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1521 = 7'h47 == _myNewVec_117_T_3[6:0] ? myVec_71 : _GEN_1520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1522 = 7'h48 == _myNewVec_117_T_3[6:0] ? myVec_72 : _GEN_1521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1523 = 7'h49 == _myNewVec_117_T_3[6:0] ? myVec_73 : _GEN_1522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1524 = 7'h4a == _myNewVec_117_T_3[6:0] ? myVec_74 : _GEN_1523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1525 = 7'h4b == _myNewVec_117_T_3[6:0] ? myVec_75 : _GEN_1524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1526 = 7'h4c == _myNewVec_117_T_3[6:0] ? myVec_76 : _GEN_1525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1527 = 7'h4d == _myNewVec_117_T_3[6:0] ? myVec_77 : _GEN_1526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1528 = 7'h4e == _myNewVec_117_T_3[6:0] ? myVec_78 : _GEN_1527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1529 = 7'h4f == _myNewVec_117_T_3[6:0] ? myVec_79 : _GEN_1528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1530 = 7'h50 == _myNewVec_117_T_3[6:0] ? myVec_80 : _GEN_1529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1531 = 7'h51 == _myNewVec_117_T_3[6:0] ? myVec_81 : _GEN_1530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1532 = 7'h52 == _myNewVec_117_T_3[6:0] ? myVec_82 : _GEN_1531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1533 = 7'h53 == _myNewVec_117_T_3[6:0] ? myVec_83 : _GEN_1532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1534 = 7'h54 == _myNewVec_117_T_3[6:0] ? myVec_84 : _GEN_1533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1535 = 7'h55 == _myNewVec_117_T_3[6:0] ? myVec_85 : _GEN_1534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1536 = 7'h56 == _myNewVec_117_T_3[6:0] ? myVec_86 : _GEN_1535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1537 = 7'h57 == _myNewVec_117_T_3[6:0] ? myVec_87 : _GEN_1536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1538 = 7'h58 == _myNewVec_117_T_3[6:0] ? myVec_88 : _GEN_1537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1539 = 7'h59 == _myNewVec_117_T_3[6:0] ? myVec_89 : _GEN_1538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1540 = 7'h5a == _myNewVec_117_T_3[6:0] ? myVec_90 : _GEN_1539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1541 = 7'h5b == _myNewVec_117_T_3[6:0] ? myVec_91 : _GEN_1540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1542 = 7'h5c == _myNewVec_117_T_3[6:0] ? myVec_92 : _GEN_1541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1543 = 7'h5d == _myNewVec_117_T_3[6:0] ? myVec_93 : _GEN_1542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1544 = 7'h5e == _myNewVec_117_T_3[6:0] ? myVec_94 : _GEN_1543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1545 = 7'h5f == _myNewVec_117_T_3[6:0] ? myVec_95 : _GEN_1544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1546 = 7'h60 == _myNewVec_117_T_3[6:0] ? myVec_96 : _GEN_1545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1547 = 7'h61 == _myNewVec_117_T_3[6:0] ? myVec_97 : _GEN_1546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1548 = 7'h62 == _myNewVec_117_T_3[6:0] ? myVec_98 : _GEN_1547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1549 = 7'h63 == _myNewVec_117_T_3[6:0] ? myVec_99 : _GEN_1548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1550 = 7'h64 == _myNewVec_117_T_3[6:0] ? myVec_100 : _GEN_1549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1551 = 7'h65 == _myNewVec_117_T_3[6:0] ? myVec_101 : _GEN_1550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1552 = 7'h66 == _myNewVec_117_T_3[6:0] ? myVec_102 : _GEN_1551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1553 = 7'h67 == _myNewVec_117_T_3[6:0] ? myVec_103 : _GEN_1552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1554 = 7'h68 == _myNewVec_117_T_3[6:0] ? myVec_104 : _GEN_1553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1555 = 7'h69 == _myNewVec_117_T_3[6:0] ? myVec_105 : _GEN_1554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1556 = 7'h6a == _myNewVec_117_T_3[6:0] ? myVec_106 : _GEN_1555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1557 = 7'h6b == _myNewVec_117_T_3[6:0] ? myVec_107 : _GEN_1556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1558 = 7'h6c == _myNewVec_117_T_3[6:0] ? myVec_108 : _GEN_1557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1559 = 7'h6d == _myNewVec_117_T_3[6:0] ? myVec_109 : _GEN_1558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1560 = 7'h6e == _myNewVec_117_T_3[6:0] ? myVec_110 : _GEN_1559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1561 = 7'h6f == _myNewVec_117_T_3[6:0] ? myVec_111 : _GEN_1560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1562 = 7'h70 == _myNewVec_117_T_3[6:0] ? myVec_112 : _GEN_1561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1563 = 7'h71 == _myNewVec_117_T_3[6:0] ? myVec_113 : _GEN_1562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1564 = 7'h72 == _myNewVec_117_T_3[6:0] ? myVec_114 : _GEN_1563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1565 = 7'h73 == _myNewVec_117_T_3[6:0] ? myVec_115 : _GEN_1564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1566 = 7'h74 == _myNewVec_117_T_3[6:0] ? myVec_116 : _GEN_1565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1567 = 7'h75 == _myNewVec_117_T_3[6:0] ? myVec_117 : _GEN_1566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1568 = 7'h76 == _myNewVec_117_T_3[6:0] ? myVec_118 : _GEN_1567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1569 = 7'h77 == _myNewVec_117_T_3[6:0] ? myVec_119 : _GEN_1568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1570 = 7'h78 == _myNewVec_117_T_3[6:0] ? myVec_120 : _GEN_1569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1571 = 7'h79 == _myNewVec_117_T_3[6:0] ? myVec_121 : _GEN_1570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1572 = 7'h7a == _myNewVec_117_T_3[6:0] ? myVec_122 : _GEN_1571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1573 = 7'h7b == _myNewVec_117_T_3[6:0] ? myVec_123 : _GEN_1572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1574 = 7'h7c == _myNewVec_117_T_3[6:0] ? myVec_124 : _GEN_1573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1575 = 7'h7d == _myNewVec_117_T_3[6:0] ? myVec_125 : _GEN_1574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1576 = 7'h7e == _myNewVec_117_T_3[6:0] ? myVec_126 : _GEN_1575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_117 = 7'h7f == _myNewVec_117_T_3[6:0] ? myVec_127 : _GEN_1576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_116_T_3 = _myNewVec_127_T_1 + 16'hb; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1579 = 7'h1 == _myNewVec_116_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1580 = 7'h2 == _myNewVec_116_T_3[6:0] ? myVec_2 : _GEN_1579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1581 = 7'h3 == _myNewVec_116_T_3[6:0] ? myVec_3 : _GEN_1580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1582 = 7'h4 == _myNewVec_116_T_3[6:0] ? myVec_4 : _GEN_1581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1583 = 7'h5 == _myNewVec_116_T_3[6:0] ? myVec_5 : _GEN_1582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1584 = 7'h6 == _myNewVec_116_T_3[6:0] ? myVec_6 : _GEN_1583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1585 = 7'h7 == _myNewVec_116_T_3[6:0] ? myVec_7 : _GEN_1584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1586 = 7'h8 == _myNewVec_116_T_3[6:0] ? myVec_8 : _GEN_1585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1587 = 7'h9 == _myNewVec_116_T_3[6:0] ? myVec_9 : _GEN_1586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1588 = 7'ha == _myNewVec_116_T_3[6:0] ? myVec_10 : _GEN_1587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1589 = 7'hb == _myNewVec_116_T_3[6:0] ? myVec_11 : _GEN_1588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1590 = 7'hc == _myNewVec_116_T_3[6:0] ? myVec_12 : _GEN_1589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1591 = 7'hd == _myNewVec_116_T_3[6:0] ? myVec_13 : _GEN_1590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1592 = 7'he == _myNewVec_116_T_3[6:0] ? myVec_14 : _GEN_1591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1593 = 7'hf == _myNewVec_116_T_3[6:0] ? myVec_15 : _GEN_1592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1594 = 7'h10 == _myNewVec_116_T_3[6:0] ? myVec_16 : _GEN_1593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1595 = 7'h11 == _myNewVec_116_T_3[6:0] ? myVec_17 : _GEN_1594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1596 = 7'h12 == _myNewVec_116_T_3[6:0] ? myVec_18 : _GEN_1595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1597 = 7'h13 == _myNewVec_116_T_3[6:0] ? myVec_19 : _GEN_1596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1598 = 7'h14 == _myNewVec_116_T_3[6:0] ? myVec_20 : _GEN_1597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1599 = 7'h15 == _myNewVec_116_T_3[6:0] ? myVec_21 : _GEN_1598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1600 = 7'h16 == _myNewVec_116_T_3[6:0] ? myVec_22 : _GEN_1599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1601 = 7'h17 == _myNewVec_116_T_3[6:0] ? myVec_23 : _GEN_1600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1602 = 7'h18 == _myNewVec_116_T_3[6:0] ? myVec_24 : _GEN_1601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1603 = 7'h19 == _myNewVec_116_T_3[6:0] ? myVec_25 : _GEN_1602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1604 = 7'h1a == _myNewVec_116_T_3[6:0] ? myVec_26 : _GEN_1603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1605 = 7'h1b == _myNewVec_116_T_3[6:0] ? myVec_27 : _GEN_1604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1606 = 7'h1c == _myNewVec_116_T_3[6:0] ? myVec_28 : _GEN_1605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1607 = 7'h1d == _myNewVec_116_T_3[6:0] ? myVec_29 : _GEN_1606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1608 = 7'h1e == _myNewVec_116_T_3[6:0] ? myVec_30 : _GEN_1607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1609 = 7'h1f == _myNewVec_116_T_3[6:0] ? myVec_31 : _GEN_1608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1610 = 7'h20 == _myNewVec_116_T_3[6:0] ? myVec_32 : _GEN_1609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1611 = 7'h21 == _myNewVec_116_T_3[6:0] ? myVec_33 : _GEN_1610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1612 = 7'h22 == _myNewVec_116_T_3[6:0] ? myVec_34 : _GEN_1611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1613 = 7'h23 == _myNewVec_116_T_3[6:0] ? myVec_35 : _GEN_1612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1614 = 7'h24 == _myNewVec_116_T_3[6:0] ? myVec_36 : _GEN_1613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1615 = 7'h25 == _myNewVec_116_T_3[6:0] ? myVec_37 : _GEN_1614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1616 = 7'h26 == _myNewVec_116_T_3[6:0] ? myVec_38 : _GEN_1615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1617 = 7'h27 == _myNewVec_116_T_3[6:0] ? myVec_39 : _GEN_1616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1618 = 7'h28 == _myNewVec_116_T_3[6:0] ? myVec_40 : _GEN_1617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1619 = 7'h29 == _myNewVec_116_T_3[6:0] ? myVec_41 : _GEN_1618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1620 = 7'h2a == _myNewVec_116_T_3[6:0] ? myVec_42 : _GEN_1619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1621 = 7'h2b == _myNewVec_116_T_3[6:0] ? myVec_43 : _GEN_1620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1622 = 7'h2c == _myNewVec_116_T_3[6:0] ? myVec_44 : _GEN_1621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1623 = 7'h2d == _myNewVec_116_T_3[6:0] ? myVec_45 : _GEN_1622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1624 = 7'h2e == _myNewVec_116_T_3[6:0] ? myVec_46 : _GEN_1623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1625 = 7'h2f == _myNewVec_116_T_3[6:0] ? myVec_47 : _GEN_1624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1626 = 7'h30 == _myNewVec_116_T_3[6:0] ? myVec_48 : _GEN_1625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1627 = 7'h31 == _myNewVec_116_T_3[6:0] ? myVec_49 : _GEN_1626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1628 = 7'h32 == _myNewVec_116_T_3[6:0] ? myVec_50 : _GEN_1627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1629 = 7'h33 == _myNewVec_116_T_3[6:0] ? myVec_51 : _GEN_1628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1630 = 7'h34 == _myNewVec_116_T_3[6:0] ? myVec_52 : _GEN_1629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1631 = 7'h35 == _myNewVec_116_T_3[6:0] ? myVec_53 : _GEN_1630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1632 = 7'h36 == _myNewVec_116_T_3[6:0] ? myVec_54 : _GEN_1631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1633 = 7'h37 == _myNewVec_116_T_3[6:0] ? myVec_55 : _GEN_1632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1634 = 7'h38 == _myNewVec_116_T_3[6:0] ? myVec_56 : _GEN_1633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1635 = 7'h39 == _myNewVec_116_T_3[6:0] ? myVec_57 : _GEN_1634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1636 = 7'h3a == _myNewVec_116_T_3[6:0] ? myVec_58 : _GEN_1635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1637 = 7'h3b == _myNewVec_116_T_3[6:0] ? myVec_59 : _GEN_1636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1638 = 7'h3c == _myNewVec_116_T_3[6:0] ? myVec_60 : _GEN_1637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1639 = 7'h3d == _myNewVec_116_T_3[6:0] ? myVec_61 : _GEN_1638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1640 = 7'h3e == _myNewVec_116_T_3[6:0] ? myVec_62 : _GEN_1639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1641 = 7'h3f == _myNewVec_116_T_3[6:0] ? myVec_63 : _GEN_1640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1642 = 7'h40 == _myNewVec_116_T_3[6:0] ? myVec_64 : _GEN_1641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1643 = 7'h41 == _myNewVec_116_T_3[6:0] ? myVec_65 : _GEN_1642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1644 = 7'h42 == _myNewVec_116_T_3[6:0] ? myVec_66 : _GEN_1643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1645 = 7'h43 == _myNewVec_116_T_3[6:0] ? myVec_67 : _GEN_1644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1646 = 7'h44 == _myNewVec_116_T_3[6:0] ? myVec_68 : _GEN_1645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1647 = 7'h45 == _myNewVec_116_T_3[6:0] ? myVec_69 : _GEN_1646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1648 = 7'h46 == _myNewVec_116_T_3[6:0] ? myVec_70 : _GEN_1647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1649 = 7'h47 == _myNewVec_116_T_3[6:0] ? myVec_71 : _GEN_1648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1650 = 7'h48 == _myNewVec_116_T_3[6:0] ? myVec_72 : _GEN_1649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1651 = 7'h49 == _myNewVec_116_T_3[6:0] ? myVec_73 : _GEN_1650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1652 = 7'h4a == _myNewVec_116_T_3[6:0] ? myVec_74 : _GEN_1651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1653 = 7'h4b == _myNewVec_116_T_3[6:0] ? myVec_75 : _GEN_1652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1654 = 7'h4c == _myNewVec_116_T_3[6:0] ? myVec_76 : _GEN_1653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1655 = 7'h4d == _myNewVec_116_T_3[6:0] ? myVec_77 : _GEN_1654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1656 = 7'h4e == _myNewVec_116_T_3[6:0] ? myVec_78 : _GEN_1655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1657 = 7'h4f == _myNewVec_116_T_3[6:0] ? myVec_79 : _GEN_1656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1658 = 7'h50 == _myNewVec_116_T_3[6:0] ? myVec_80 : _GEN_1657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1659 = 7'h51 == _myNewVec_116_T_3[6:0] ? myVec_81 : _GEN_1658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1660 = 7'h52 == _myNewVec_116_T_3[6:0] ? myVec_82 : _GEN_1659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1661 = 7'h53 == _myNewVec_116_T_3[6:0] ? myVec_83 : _GEN_1660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1662 = 7'h54 == _myNewVec_116_T_3[6:0] ? myVec_84 : _GEN_1661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1663 = 7'h55 == _myNewVec_116_T_3[6:0] ? myVec_85 : _GEN_1662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1664 = 7'h56 == _myNewVec_116_T_3[6:0] ? myVec_86 : _GEN_1663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1665 = 7'h57 == _myNewVec_116_T_3[6:0] ? myVec_87 : _GEN_1664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1666 = 7'h58 == _myNewVec_116_T_3[6:0] ? myVec_88 : _GEN_1665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1667 = 7'h59 == _myNewVec_116_T_3[6:0] ? myVec_89 : _GEN_1666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1668 = 7'h5a == _myNewVec_116_T_3[6:0] ? myVec_90 : _GEN_1667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1669 = 7'h5b == _myNewVec_116_T_3[6:0] ? myVec_91 : _GEN_1668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1670 = 7'h5c == _myNewVec_116_T_3[6:0] ? myVec_92 : _GEN_1669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1671 = 7'h5d == _myNewVec_116_T_3[6:0] ? myVec_93 : _GEN_1670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1672 = 7'h5e == _myNewVec_116_T_3[6:0] ? myVec_94 : _GEN_1671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1673 = 7'h5f == _myNewVec_116_T_3[6:0] ? myVec_95 : _GEN_1672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1674 = 7'h60 == _myNewVec_116_T_3[6:0] ? myVec_96 : _GEN_1673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1675 = 7'h61 == _myNewVec_116_T_3[6:0] ? myVec_97 : _GEN_1674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1676 = 7'h62 == _myNewVec_116_T_3[6:0] ? myVec_98 : _GEN_1675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1677 = 7'h63 == _myNewVec_116_T_3[6:0] ? myVec_99 : _GEN_1676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1678 = 7'h64 == _myNewVec_116_T_3[6:0] ? myVec_100 : _GEN_1677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1679 = 7'h65 == _myNewVec_116_T_3[6:0] ? myVec_101 : _GEN_1678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1680 = 7'h66 == _myNewVec_116_T_3[6:0] ? myVec_102 : _GEN_1679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1681 = 7'h67 == _myNewVec_116_T_3[6:0] ? myVec_103 : _GEN_1680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1682 = 7'h68 == _myNewVec_116_T_3[6:0] ? myVec_104 : _GEN_1681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1683 = 7'h69 == _myNewVec_116_T_3[6:0] ? myVec_105 : _GEN_1682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1684 = 7'h6a == _myNewVec_116_T_3[6:0] ? myVec_106 : _GEN_1683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1685 = 7'h6b == _myNewVec_116_T_3[6:0] ? myVec_107 : _GEN_1684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1686 = 7'h6c == _myNewVec_116_T_3[6:0] ? myVec_108 : _GEN_1685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1687 = 7'h6d == _myNewVec_116_T_3[6:0] ? myVec_109 : _GEN_1686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1688 = 7'h6e == _myNewVec_116_T_3[6:0] ? myVec_110 : _GEN_1687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1689 = 7'h6f == _myNewVec_116_T_3[6:0] ? myVec_111 : _GEN_1688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1690 = 7'h70 == _myNewVec_116_T_3[6:0] ? myVec_112 : _GEN_1689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1691 = 7'h71 == _myNewVec_116_T_3[6:0] ? myVec_113 : _GEN_1690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1692 = 7'h72 == _myNewVec_116_T_3[6:0] ? myVec_114 : _GEN_1691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1693 = 7'h73 == _myNewVec_116_T_3[6:0] ? myVec_115 : _GEN_1692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1694 = 7'h74 == _myNewVec_116_T_3[6:0] ? myVec_116 : _GEN_1693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1695 = 7'h75 == _myNewVec_116_T_3[6:0] ? myVec_117 : _GEN_1694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1696 = 7'h76 == _myNewVec_116_T_3[6:0] ? myVec_118 : _GEN_1695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1697 = 7'h77 == _myNewVec_116_T_3[6:0] ? myVec_119 : _GEN_1696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1698 = 7'h78 == _myNewVec_116_T_3[6:0] ? myVec_120 : _GEN_1697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1699 = 7'h79 == _myNewVec_116_T_3[6:0] ? myVec_121 : _GEN_1698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1700 = 7'h7a == _myNewVec_116_T_3[6:0] ? myVec_122 : _GEN_1699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1701 = 7'h7b == _myNewVec_116_T_3[6:0] ? myVec_123 : _GEN_1700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1702 = 7'h7c == _myNewVec_116_T_3[6:0] ? myVec_124 : _GEN_1701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1703 = 7'h7d == _myNewVec_116_T_3[6:0] ? myVec_125 : _GEN_1702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1704 = 7'h7e == _myNewVec_116_T_3[6:0] ? myVec_126 : _GEN_1703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_116 = 7'h7f == _myNewVec_116_T_3[6:0] ? myVec_127 : _GEN_1704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_115_T_3 = _myNewVec_127_T_1 + 16'hc; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1707 = 7'h1 == _myNewVec_115_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1708 = 7'h2 == _myNewVec_115_T_3[6:0] ? myVec_2 : _GEN_1707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1709 = 7'h3 == _myNewVec_115_T_3[6:0] ? myVec_3 : _GEN_1708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1710 = 7'h4 == _myNewVec_115_T_3[6:0] ? myVec_4 : _GEN_1709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1711 = 7'h5 == _myNewVec_115_T_3[6:0] ? myVec_5 : _GEN_1710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1712 = 7'h6 == _myNewVec_115_T_3[6:0] ? myVec_6 : _GEN_1711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1713 = 7'h7 == _myNewVec_115_T_3[6:0] ? myVec_7 : _GEN_1712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1714 = 7'h8 == _myNewVec_115_T_3[6:0] ? myVec_8 : _GEN_1713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1715 = 7'h9 == _myNewVec_115_T_3[6:0] ? myVec_9 : _GEN_1714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1716 = 7'ha == _myNewVec_115_T_3[6:0] ? myVec_10 : _GEN_1715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1717 = 7'hb == _myNewVec_115_T_3[6:0] ? myVec_11 : _GEN_1716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1718 = 7'hc == _myNewVec_115_T_3[6:0] ? myVec_12 : _GEN_1717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1719 = 7'hd == _myNewVec_115_T_3[6:0] ? myVec_13 : _GEN_1718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1720 = 7'he == _myNewVec_115_T_3[6:0] ? myVec_14 : _GEN_1719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1721 = 7'hf == _myNewVec_115_T_3[6:0] ? myVec_15 : _GEN_1720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1722 = 7'h10 == _myNewVec_115_T_3[6:0] ? myVec_16 : _GEN_1721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1723 = 7'h11 == _myNewVec_115_T_3[6:0] ? myVec_17 : _GEN_1722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1724 = 7'h12 == _myNewVec_115_T_3[6:0] ? myVec_18 : _GEN_1723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1725 = 7'h13 == _myNewVec_115_T_3[6:0] ? myVec_19 : _GEN_1724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1726 = 7'h14 == _myNewVec_115_T_3[6:0] ? myVec_20 : _GEN_1725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1727 = 7'h15 == _myNewVec_115_T_3[6:0] ? myVec_21 : _GEN_1726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1728 = 7'h16 == _myNewVec_115_T_3[6:0] ? myVec_22 : _GEN_1727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1729 = 7'h17 == _myNewVec_115_T_3[6:0] ? myVec_23 : _GEN_1728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1730 = 7'h18 == _myNewVec_115_T_3[6:0] ? myVec_24 : _GEN_1729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1731 = 7'h19 == _myNewVec_115_T_3[6:0] ? myVec_25 : _GEN_1730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1732 = 7'h1a == _myNewVec_115_T_3[6:0] ? myVec_26 : _GEN_1731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1733 = 7'h1b == _myNewVec_115_T_3[6:0] ? myVec_27 : _GEN_1732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1734 = 7'h1c == _myNewVec_115_T_3[6:0] ? myVec_28 : _GEN_1733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1735 = 7'h1d == _myNewVec_115_T_3[6:0] ? myVec_29 : _GEN_1734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1736 = 7'h1e == _myNewVec_115_T_3[6:0] ? myVec_30 : _GEN_1735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1737 = 7'h1f == _myNewVec_115_T_3[6:0] ? myVec_31 : _GEN_1736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1738 = 7'h20 == _myNewVec_115_T_3[6:0] ? myVec_32 : _GEN_1737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1739 = 7'h21 == _myNewVec_115_T_3[6:0] ? myVec_33 : _GEN_1738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1740 = 7'h22 == _myNewVec_115_T_3[6:0] ? myVec_34 : _GEN_1739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1741 = 7'h23 == _myNewVec_115_T_3[6:0] ? myVec_35 : _GEN_1740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1742 = 7'h24 == _myNewVec_115_T_3[6:0] ? myVec_36 : _GEN_1741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1743 = 7'h25 == _myNewVec_115_T_3[6:0] ? myVec_37 : _GEN_1742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1744 = 7'h26 == _myNewVec_115_T_3[6:0] ? myVec_38 : _GEN_1743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1745 = 7'h27 == _myNewVec_115_T_3[6:0] ? myVec_39 : _GEN_1744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1746 = 7'h28 == _myNewVec_115_T_3[6:0] ? myVec_40 : _GEN_1745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1747 = 7'h29 == _myNewVec_115_T_3[6:0] ? myVec_41 : _GEN_1746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1748 = 7'h2a == _myNewVec_115_T_3[6:0] ? myVec_42 : _GEN_1747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1749 = 7'h2b == _myNewVec_115_T_3[6:0] ? myVec_43 : _GEN_1748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1750 = 7'h2c == _myNewVec_115_T_3[6:0] ? myVec_44 : _GEN_1749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1751 = 7'h2d == _myNewVec_115_T_3[6:0] ? myVec_45 : _GEN_1750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1752 = 7'h2e == _myNewVec_115_T_3[6:0] ? myVec_46 : _GEN_1751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1753 = 7'h2f == _myNewVec_115_T_3[6:0] ? myVec_47 : _GEN_1752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1754 = 7'h30 == _myNewVec_115_T_3[6:0] ? myVec_48 : _GEN_1753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1755 = 7'h31 == _myNewVec_115_T_3[6:0] ? myVec_49 : _GEN_1754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1756 = 7'h32 == _myNewVec_115_T_3[6:0] ? myVec_50 : _GEN_1755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1757 = 7'h33 == _myNewVec_115_T_3[6:0] ? myVec_51 : _GEN_1756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1758 = 7'h34 == _myNewVec_115_T_3[6:0] ? myVec_52 : _GEN_1757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1759 = 7'h35 == _myNewVec_115_T_3[6:0] ? myVec_53 : _GEN_1758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1760 = 7'h36 == _myNewVec_115_T_3[6:0] ? myVec_54 : _GEN_1759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1761 = 7'h37 == _myNewVec_115_T_3[6:0] ? myVec_55 : _GEN_1760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1762 = 7'h38 == _myNewVec_115_T_3[6:0] ? myVec_56 : _GEN_1761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1763 = 7'h39 == _myNewVec_115_T_3[6:0] ? myVec_57 : _GEN_1762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1764 = 7'h3a == _myNewVec_115_T_3[6:0] ? myVec_58 : _GEN_1763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1765 = 7'h3b == _myNewVec_115_T_3[6:0] ? myVec_59 : _GEN_1764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1766 = 7'h3c == _myNewVec_115_T_3[6:0] ? myVec_60 : _GEN_1765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1767 = 7'h3d == _myNewVec_115_T_3[6:0] ? myVec_61 : _GEN_1766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1768 = 7'h3e == _myNewVec_115_T_3[6:0] ? myVec_62 : _GEN_1767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1769 = 7'h3f == _myNewVec_115_T_3[6:0] ? myVec_63 : _GEN_1768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1770 = 7'h40 == _myNewVec_115_T_3[6:0] ? myVec_64 : _GEN_1769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1771 = 7'h41 == _myNewVec_115_T_3[6:0] ? myVec_65 : _GEN_1770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1772 = 7'h42 == _myNewVec_115_T_3[6:0] ? myVec_66 : _GEN_1771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1773 = 7'h43 == _myNewVec_115_T_3[6:0] ? myVec_67 : _GEN_1772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1774 = 7'h44 == _myNewVec_115_T_3[6:0] ? myVec_68 : _GEN_1773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1775 = 7'h45 == _myNewVec_115_T_3[6:0] ? myVec_69 : _GEN_1774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1776 = 7'h46 == _myNewVec_115_T_3[6:0] ? myVec_70 : _GEN_1775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1777 = 7'h47 == _myNewVec_115_T_3[6:0] ? myVec_71 : _GEN_1776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1778 = 7'h48 == _myNewVec_115_T_3[6:0] ? myVec_72 : _GEN_1777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1779 = 7'h49 == _myNewVec_115_T_3[6:0] ? myVec_73 : _GEN_1778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1780 = 7'h4a == _myNewVec_115_T_3[6:0] ? myVec_74 : _GEN_1779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1781 = 7'h4b == _myNewVec_115_T_3[6:0] ? myVec_75 : _GEN_1780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1782 = 7'h4c == _myNewVec_115_T_3[6:0] ? myVec_76 : _GEN_1781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1783 = 7'h4d == _myNewVec_115_T_3[6:0] ? myVec_77 : _GEN_1782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1784 = 7'h4e == _myNewVec_115_T_3[6:0] ? myVec_78 : _GEN_1783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1785 = 7'h4f == _myNewVec_115_T_3[6:0] ? myVec_79 : _GEN_1784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1786 = 7'h50 == _myNewVec_115_T_3[6:0] ? myVec_80 : _GEN_1785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1787 = 7'h51 == _myNewVec_115_T_3[6:0] ? myVec_81 : _GEN_1786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1788 = 7'h52 == _myNewVec_115_T_3[6:0] ? myVec_82 : _GEN_1787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1789 = 7'h53 == _myNewVec_115_T_3[6:0] ? myVec_83 : _GEN_1788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1790 = 7'h54 == _myNewVec_115_T_3[6:0] ? myVec_84 : _GEN_1789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1791 = 7'h55 == _myNewVec_115_T_3[6:0] ? myVec_85 : _GEN_1790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1792 = 7'h56 == _myNewVec_115_T_3[6:0] ? myVec_86 : _GEN_1791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1793 = 7'h57 == _myNewVec_115_T_3[6:0] ? myVec_87 : _GEN_1792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1794 = 7'h58 == _myNewVec_115_T_3[6:0] ? myVec_88 : _GEN_1793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1795 = 7'h59 == _myNewVec_115_T_3[6:0] ? myVec_89 : _GEN_1794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1796 = 7'h5a == _myNewVec_115_T_3[6:0] ? myVec_90 : _GEN_1795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1797 = 7'h5b == _myNewVec_115_T_3[6:0] ? myVec_91 : _GEN_1796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1798 = 7'h5c == _myNewVec_115_T_3[6:0] ? myVec_92 : _GEN_1797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1799 = 7'h5d == _myNewVec_115_T_3[6:0] ? myVec_93 : _GEN_1798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1800 = 7'h5e == _myNewVec_115_T_3[6:0] ? myVec_94 : _GEN_1799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1801 = 7'h5f == _myNewVec_115_T_3[6:0] ? myVec_95 : _GEN_1800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1802 = 7'h60 == _myNewVec_115_T_3[6:0] ? myVec_96 : _GEN_1801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1803 = 7'h61 == _myNewVec_115_T_3[6:0] ? myVec_97 : _GEN_1802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1804 = 7'h62 == _myNewVec_115_T_3[6:0] ? myVec_98 : _GEN_1803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1805 = 7'h63 == _myNewVec_115_T_3[6:0] ? myVec_99 : _GEN_1804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1806 = 7'h64 == _myNewVec_115_T_3[6:0] ? myVec_100 : _GEN_1805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1807 = 7'h65 == _myNewVec_115_T_3[6:0] ? myVec_101 : _GEN_1806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1808 = 7'h66 == _myNewVec_115_T_3[6:0] ? myVec_102 : _GEN_1807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1809 = 7'h67 == _myNewVec_115_T_3[6:0] ? myVec_103 : _GEN_1808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1810 = 7'h68 == _myNewVec_115_T_3[6:0] ? myVec_104 : _GEN_1809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1811 = 7'h69 == _myNewVec_115_T_3[6:0] ? myVec_105 : _GEN_1810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1812 = 7'h6a == _myNewVec_115_T_3[6:0] ? myVec_106 : _GEN_1811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1813 = 7'h6b == _myNewVec_115_T_3[6:0] ? myVec_107 : _GEN_1812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1814 = 7'h6c == _myNewVec_115_T_3[6:0] ? myVec_108 : _GEN_1813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1815 = 7'h6d == _myNewVec_115_T_3[6:0] ? myVec_109 : _GEN_1814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1816 = 7'h6e == _myNewVec_115_T_3[6:0] ? myVec_110 : _GEN_1815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1817 = 7'h6f == _myNewVec_115_T_3[6:0] ? myVec_111 : _GEN_1816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1818 = 7'h70 == _myNewVec_115_T_3[6:0] ? myVec_112 : _GEN_1817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1819 = 7'h71 == _myNewVec_115_T_3[6:0] ? myVec_113 : _GEN_1818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1820 = 7'h72 == _myNewVec_115_T_3[6:0] ? myVec_114 : _GEN_1819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1821 = 7'h73 == _myNewVec_115_T_3[6:0] ? myVec_115 : _GEN_1820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1822 = 7'h74 == _myNewVec_115_T_3[6:0] ? myVec_116 : _GEN_1821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1823 = 7'h75 == _myNewVec_115_T_3[6:0] ? myVec_117 : _GEN_1822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1824 = 7'h76 == _myNewVec_115_T_3[6:0] ? myVec_118 : _GEN_1823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1825 = 7'h77 == _myNewVec_115_T_3[6:0] ? myVec_119 : _GEN_1824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1826 = 7'h78 == _myNewVec_115_T_3[6:0] ? myVec_120 : _GEN_1825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1827 = 7'h79 == _myNewVec_115_T_3[6:0] ? myVec_121 : _GEN_1826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1828 = 7'h7a == _myNewVec_115_T_3[6:0] ? myVec_122 : _GEN_1827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1829 = 7'h7b == _myNewVec_115_T_3[6:0] ? myVec_123 : _GEN_1828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1830 = 7'h7c == _myNewVec_115_T_3[6:0] ? myVec_124 : _GEN_1829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1831 = 7'h7d == _myNewVec_115_T_3[6:0] ? myVec_125 : _GEN_1830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1832 = 7'h7e == _myNewVec_115_T_3[6:0] ? myVec_126 : _GEN_1831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_115 = 7'h7f == _myNewVec_115_T_3[6:0] ? myVec_127 : _GEN_1832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_114_T_3 = _myNewVec_127_T_1 + 16'hd; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1835 = 7'h1 == _myNewVec_114_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1836 = 7'h2 == _myNewVec_114_T_3[6:0] ? myVec_2 : _GEN_1835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1837 = 7'h3 == _myNewVec_114_T_3[6:0] ? myVec_3 : _GEN_1836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1838 = 7'h4 == _myNewVec_114_T_3[6:0] ? myVec_4 : _GEN_1837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1839 = 7'h5 == _myNewVec_114_T_3[6:0] ? myVec_5 : _GEN_1838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1840 = 7'h6 == _myNewVec_114_T_3[6:0] ? myVec_6 : _GEN_1839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1841 = 7'h7 == _myNewVec_114_T_3[6:0] ? myVec_7 : _GEN_1840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1842 = 7'h8 == _myNewVec_114_T_3[6:0] ? myVec_8 : _GEN_1841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1843 = 7'h9 == _myNewVec_114_T_3[6:0] ? myVec_9 : _GEN_1842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1844 = 7'ha == _myNewVec_114_T_3[6:0] ? myVec_10 : _GEN_1843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1845 = 7'hb == _myNewVec_114_T_3[6:0] ? myVec_11 : _GEN_1844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1846 = 7'hc == _myNewVec_114_T_3[6:0] ? myVec_12 : _GEN_1845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1847 = 7'hd == _myNewVec_114_T_3[6:0] ? myVec_13 : _GEN_1846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1848 = 7'he == _myNewVec_114_T_3[6:0] ? myVec_14 : _GEN_1847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1849 = 7'hf == _myNewVec_114_T_3[6:0] ? myVec_15 : _GEN_1848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1850 = 7'h10 == _myNewVec_114_T_3[6:0] ? myVec_16 : _GEN_1849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1851 = 7'h11 == _myNewVec_114_T_3[6:0] ? myVec_17 : _GEN_1850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1852 = 7'h12 == _myNewVec_114_T_3[6:0] ? myVec_18 : _GEN_1851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1853 = 7'h13 == _myNewVec_114_T_3[6:0] ? myVec_19 : _GEN_1852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1854 = 7'h14 == _myNewVec_114_T_3[6:0] ? myVec_20 : _GEN_1853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1855 = 7'h15 == _myNewVec_114_T_3[6:0] ? myVec_21 : _GEN_1854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1856 = 7'h16 == _myNewVec_114_T_3[6:0] ? myVec_22 : _GEN_1855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1857 = 7'h17 == _myNewVec_114_T_3[6:0] ? myVec_23 : _GEN_1856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1858 = 7'h18 == _myNewVec_114_T_3[6:0] ? myVec_24 : _GEN_1857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1859 = 7'h19 == _myNewVec_114_T_3[6:0] ? myVec_25 : _GEN_1858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1860 = 7'h1a == _myNewVec_114_T_3[6:0] ? myVec_26 : _GEN_1859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1861 = 7'h1b == _myNewVec_114_T_3[6:0] ? myVec_27 : _GEN_1860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1862 = 7'h1c == _myNewVec_114_T_3[6:0] ? myVec_28 : _GEN_1861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1863 = 7'h1d == _myNewVec_114_T_3[6:0] ? myVec_29 : _GEN_1862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1864 = 7'h1e == _myNewVec_114_T_3[6:0] ? myVec_30 : _GEN_1863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1865 = 7'h1f == _myNewVec_114_T_3[6:0] ? myVec_31 : _GEN_1864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1866 = 7'h20 == _myNewVec_114_T_3[6:0] ? myVec_32 : _GEN_1865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1867 = 7'h21 == _myNewVec_114_T_3[6:0] ? myVec_33 : _GEN_1866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1868 = 7'h22 == _myNewVec_114_T_3[6:0] ? myVec_34 : _GEN_1867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1869 = 7'h23 == _myNewVec_114_T_3[6:0] ? myVec_35 : _GEN_1868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1870 = 7'h24 == _myNewVec_114_T_3[6:0] ? myVec_36 : _GEN_1869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1871 = 7'h25 == _myNewVec_114_T_3[6:0] ? myVec_37 : _GEN_1870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1872 = 7'h26 == _myNewVec_114_T_3[6:0] ? myVec_38 : _GEN_1871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1873 = 7'h27 == _myNewVec_114_T_3[6:0] ? myVec_39 : _GEN_1872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1874 = 7'h28 == _myNewVec_114_T_3[6:0] ? myVec_40 : _GEN_1873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1875 = 7'h29 == _myNewVec_114_T_3[6:0] ? myVec_41 : _GEN_1874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1876 = 7'h2a == _myNewVec_114_T_3[6:0] ? myVec_42 : _GEN_1875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1877 = 7'h2b == _myNewVec_114_T_3[6:0] ? myVec_43 : _GEN_1876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1878 = 7'h2c == _myNewVec_114_T_3[6:0] ? myVec_44 : _GEN_1877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1879 = 7'h2d == _myNewVec_114_T_3[6:0] ? myVec_45 : _GEN_1878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1880 = 7'h2e == _myNewVec_114_T_3[6:0] ? myVec_46 : _GEN_1879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1881 = 7'h2f == _myNewVec_114_T_3[6:0] ? myVec_47 : _GEN_1880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1882 = 7'h30 == _myNewVec_114_T_3[6:0] ? myVec_48 : _GEN_1881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1883 = 7'h31 == _myNewVec_114_T_3[6:0] ? myVec_49 : _GEN_1882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1884 = 7'h32 == _myNewVec_114_T_3[6:0] ? myVec_50 : _GEN_1883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1885 = 7'h33 == _myNewVec_114_T_3[6:0] ? myVec_51 : _GEN_1884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1886 = 7'h34 == _myNewVec_114_T_3[6:0] ? myVec_52 : _GEN_1885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1887 = 7'h35 == _myNewVec_114_T_3[6:0] ? myVec_53 : _GEN_1886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1888 = 7'h36 == _myNewVec_114_T_3[6:0] ? myVec_54 : _GEN_1887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1889 = 7'h37 == _myNewVec_114_T_3[6:0] ? myVec_55 : _GEN_1888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1890 = 7'h38 == _myNewVec_114_T_3[6:0] ? myVec_56 : _GEN_1889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1891 = 7'h39 == _myNewVec_114_T_3[6:0] ? myVec_57 : _GEN_1890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1892 = 7'h3a == _myNewVec_114_T_3[6:0] ? myVec_58 : _GEN_1891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1893 = 7'h3b == _myNewVec_114_T_3[6:0] ? myVec_59 : _GEN_1892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1894 = 7'h3c == _myNewVec_114_T_3[6:0] ? myVec_60 : _GEN_1893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1895 = 7'h3d == _myNewVec_114_T_3[6:0] ? myVec_61 : _GEN_1894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1896 = 7'h3e == _myNewVec_114_T_3[6:0] ? myVec_62 : _GEN_1895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1897 = 7'h3f == _myNewVec_114_T_3[6:0] ? myVec_63 : _GEN_1896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1898 = 7'h40 == _myNewVec_114_T_3[6:0] ? myVec_64 : _GEN_1897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1899 = 7'h41 == _myNewVec_114_T_3[6:0] ? myVec_65 : _GEN_1898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1900 = 7'h42 == _myNewVec_114_T_3[6:0] ? myVec_66 : _GEN_1899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1901 = 7'h43 == _myNewVec_114_T_3[6:0] ? myVec_67 : _GEN_1900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1902 = 7'h44 == _myNewVec_114_T_3[6:0] ? myVec_68 : _GEN_1901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1903 = 7'h45 == _myNewVec_114_T_3[6:0] ? myVec_69 : _GEN_1902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1904 = 7'h46 == _myNewVec_114_T_3[6:0] ? myVec_70 : _GEN_1903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1905 = 7'h47 == _myNewVec_114_T_3[6:0] ? myVec_71 : _GEN_1904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1906 = 7'h48 == _myNewVec_114_T_3[6:0] ? myVec_72 : _GEN_1905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1907 = 7'h49 == _myNewVec_114_T_3[6:0] ? myVec_73 : _GEN_1906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1908 = 7'h4a == _myNewVec_114_T_3[6:0] ? myVec_74 : _GEN_1907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1909 = 7'h4b == _myNewVec_114_T_3[6:0] ? myVec_75 : _GEN_1908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1910 = 7'h4c == _myNewVec_114_T_3[6:0] ? myVec_76 : _GEN_1909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1911 = 7'h4d == _myNewVec_114_T_3[6:0] ? myVec_77 : _GEN_1910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1912 = 7'h4e == _myNewVec_114_T_3[6:0] ? myVec_78 : _GEN_1911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1913 = 7'h4f == _myNewVec_114_T_3[6:0] ? myVec_79 : _GEN_1912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1914 = 7'h50 == _myNewVec_114_T_3[6:0] ? myVec_80 : _GEN_1913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1915 = 7'h51 == _myNewVec_114_T_3[6:0] ? myVec_81 : _GEN_1914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1916 = 7'h52 == _myNewVec_114_T_3[6:0] ? myVec_82 : _GEN_1915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1917 = 7'h53 == _myNewVec_114_T_3[6:0] ? myVec_83 : _GEN_1916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1918 = 7'h54 == _myNewVec_114_T_3[6:0] ? myVec_84 : _GEN_1917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1919 = 7'h55 == _myNewVec_114_T_3[6:0] ? myVec_85 : _GEN_1918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1920 = 7'h56 == _myNewVec_114_T_3[6:0] ? myVec_86 : _GEN_1919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1921 = 7'h57 == _myNewVec_114_T_3[6:0] ? myVec_87 : _GEN_1920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1922 = 7'h58 == _myNewVec_114_T_3[6:0] ? myVec_88 : _GEN_1921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1923 = 7'h59 == _myNewVec_114_T_3[6:0] ? myVec_89 : _GEN_1922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1924 = 7'h5a == _myNewVec_114_T_3[6:0] ? myVec_90 : _GEN_1923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1925 = 7'h5b == _myNewVec_114_T_3[6:0] ? myVec_91 : _GEN_1924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1926 = 7'h5c == _myNewVec_114_T_3[6:0] ? myVec_92 : _GEN_1925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1927 = 7'h5d == _myNewVec_114_T_3[6:0] ? myVec_93 : _GEN_1926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1928 = 7'h5e == _myNewVec_114_T_3[6:0] ? myVec_94 : _GEN_1927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1929 = 7'h5f == _myNewVec_114_T_3[6:0] ? myVec_95 : _GEN_1928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1930 = 7'h60 == _myNewVec_114_T_3[6:0] ? myVec_96 : _GEN_1929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1931 = 7'h61 == _myNewVec_114_T_3[6:0] ? myVec_97 : _GEN_1930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1932 = 7'h62 == _myNewVec_114_T_3[6:0] ? myVec_98 : _GEN_1931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1933 = 7'h63 == _myNewVec_114_T_3[6:0] ? myVec_99 : _GEN_1932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1934 = 7'h64 == _myNewVec_114_T_3[6:0] ? myVec_100 : _GEN_1933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1935 = 7'h65 == _myNewVec_114_T_3[6:0] ? myVec_101 : _GEN_1934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1936 = 7'h66 == _myNewVec_114_T_3[6:0] ? myVec_102 : _GEN_1935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1937 = 7'h67 == _myNewVec_114_T_3[6:0] ? myVec_103 : _GEN_1936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1938 = 7'h68 == _myNewVec_114_T_3[6:0] ? myVec_104 : _GEN_1937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1939 = 7'h69 == _myNewVec_114_T_3[6:0] ? myVec_105 : _GEN_1938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1940 = 7'h6a == _myNewVec_114_T_3[6:0] ? myVec_106 : _GEN_1939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1941 = 7'h6b == _myNewVec_114_T_3[6:0] ? myVec_107 : _GEN_1940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1942 = 7'h6c == _myNewVec_114_T_3[6:0] ? myVec_108 : _GEN_1941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1943 = 7'h6d == _myNewVec_114_T_3[6:0] ? myVec_109 : _GEN_1942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1944 = 7'h6e == _myNewVec_114_T_3[6:0] ? myVec_110 : _GEN_1943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1945 = 7'h6f == _myNewVec_114_T_3[6:0] ? myVec_111 : _GEN_1944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1946 = 7'h70 == _myNewVec_114_T_3[6:0] ? myVec_112 : _GEN_1945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1947 = 7'h71 == _myNewVec_114_T_3[6:0] ? myVec_113 : _GEN_1946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1948 = 7'h72 == _myNewVec_114_T_3[6:0] ? myVec_114 : _GEN_1947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1949 = 7'h73 == _myNewVec_114_T_3[6:0] ? myVec_115 : _GEN_1948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1950 = 7'h74 == _myNewVec_114_T_3[6:0] ? myVec_116 : _GEN_1949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1951 = 7'h75 == _myNewVec_114_T_3[6:0] ? myVec_117 : _GEN_1950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1952 = 7'h76 == _myNewVec_114_T_3[6:0] ? myVec_118 : _GEN_1951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1953 = 7'h77 == _myNewVec_114_T_3[6:0] ? myVec_119 : _GEN_1952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1954 = 7'h78 == _myNewVec_114_T_3[6:0] ? myVec_120 : _GEN_1953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1955 = 7'h79 == _myNewVec_114_T_3[6:0] ? myVec_121 : _GEN_1954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1956 = 7'h7a == _myNewVec_114_T_3[6:0] ? myVec_122 : _GEN_1955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1957 = 7'h7b == _myNewVec_114_T_3[6:0] ? myVec_123 : _GEN_1956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1958 = 7'h7c == _myNewVec_114_T_3[6:0] ? myVec_124 : _GEN_1957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1959 = 7'h7d == _myNewVec_114_T_3[6:0] ? myVec_125 : _GEN_1958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1960 = 7'h7e == _myNewVec_114_T_3[6:0] ? myVec_126 : _GEN_1959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_114 = 7'h7f == _myNewVec_114_T_3[6:0] ? myVec_127 : _GEN_1960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_113_T_3 = _myNewVec_127_T_1 + 16'he; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1963 = 7'h1 == _myNewVec_113_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1964 = 7'h2 == _myNewVec_113_T_3[6:0] ? myVec_2 : _GEN_1963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1965 = 7'h3 == _myNewVec_113_T_3[6:0] ? myVec_3 : _GEN_1964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1966 = 7'h4 == _myNewVec_113_T_3[6:0] ? myVec_4 : _GEN_1965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1967 = 7'h5 == _myNewVec_113_T_3[6:0] ? myVec_5 : _GEN_1966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1968 = 7'h6 == _myNewVec_113_T_3[6:0] ? myVec_6 : _GEN_1967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1969 = 7'h7 == _myNewVec_113_T_3[6:0] ? myVec_7 : _GEN_1968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1970 = 7'h8 == _myNewVec_113_T_3[6:0] ? myVec_8 : _GEN_1969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1971 = 7'h9 == _myNewVec_113_T_3[6:0] ? myVec_9 : _GEN_1970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1972 = 7'ha == _myNewVec_113_T_3[6:0] ? myVec_10 : _GEN_1971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1973 = 7'hb == _myNewVec_113_T_3[6:0] ? myVec_11 : _GEN_1972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1974 = 7'hc == _myNewVec_113_T_3[6:0] ? myVec_12 : _GEN_1973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1975 = 7'hd == _myNewVec_113_T_3[6:0] ? myVec_13 : _GEN_1974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1976 = 7'he == _myNewVec_113_T_3[6:0] ? myVec_14 : _GEN_1975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1977 = 7'hf == _myNewVec_113_T_3[6:0] ? myVec_15 : _GEN_1976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1978 = 7'h10 == _myNewVec_113_T_3[6:0] ? myVec_16 : _GEN_1977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1979 = 7'h11 == _myNewVec_113_T_3[6:0] ? myVec_17 : _GEN_1978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1980 = 7'h12 == _myNewVec_113_T_3[6:0] ? myVec_18 : _GEN_1979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1981 = 7'h13 == _myNewVec_113_T_3[6:0] ? myVec_19 : _GEN_1980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1982 = 7'h14 == _myNewVec_113_T_3[6:0] ? myVec_20 : _GEN_1981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1983 = 7'h15 == _myNewVec_113_T_3[6:0] ? myVec_21 : _GEN_1982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1984 = 7'h16 == _myNewVec_113_T_3[6:0] ? myVec_22 : _GEN_1983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1985 = 7'h17 == _myNewVec_113_T_3[6:0] ? myVec_23 : _GEN_1984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1986 = 7'h18 == _myNewVec_113_T_3[6:0] ? myVec_24 : _GEN_1985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1987 = 7'h19 == _myNewVec_113_T_3[6:0] ? myVec_25 : _GEN_1986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1988 = 7'h1a == _myNewVec_113_T_3[6:0] ? myVec_26 : _GEN_1987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1989 = 7'h1b == _myNewVec_113_T_3[6:0] ? myVec_27 : _GEN_1988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1990 = 7'h1c == _myNewVec_113_T_3[6:0] ? myVec_28 : _GEN_1989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1991 = 7'h1d == _myNewVec_113_T_3[6:0] ? myVec_29 : _GEN_1990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1992 = 7'h1e == _myNewVec_113_T_3[6:0] ? myVec_30 : _GEN_1991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1993 = 7'h1f == _myNewVec_113_T_3[6:0] ? myVec_31 : _GEN_1992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1994 = 7'h20 == _myNewVec_113_T_3[6:0] ? myVec_32 : _GEN_1993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1995 = 7'h21 == _myNewVec_113_T_3[6:0] ? myVec_33 : _GEN_1994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1996 = 7'h22 == _myNewVec_113_T_3[6:0] ? myVec_34 : _GEN_1995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1997 = 7'h23 == _myNewVec_113_T_3[6:0] ? myVec_35 : _GEN_1996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1998 = 7'h24 == _myNewVec_113_T_3[6:0] ? myVec_36 : _GEN_1997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1999 = 7'h25 == _myNewVec_113_T_3[6:0] ? myVec_37 : _GEN_1998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2000 = 7'h26 == _myNewVec_113_T_3[6:0] ? myVec_38 : _GEN_1999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2001 = 7'h27 == _myNewVec_113_T_3[6:0] ? myVec_39 : _GEN_2000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2002 = 7'h28 == _myNewVec_113_T_3[6:0] ? myVec_40 : _GEN_2001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2003 = 7'h29 == _myNewVec_113_T_3[6:0] ? myVec_41 : _GEN_2002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2004 = 7'h2a == _myNewVec_113_T_3[6:0] ? myVec_42 : _GEN_2003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2005 = 7'h2b == _myNewVec_113_T_3[6:0] ? myVec_43 : _GEN_2004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2006 = 7'h2c == _myNewVec_113_T_3[6:0] ? myVec_44 : _GEN_2005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2007 = 7'h2d == _myNewVec_113_T_3[6:0] ? myVec_45 : _GEN_2006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2008 = 7'h2e == _myNewVec_113_T_3[6:0] ? myVec_46 : _GEN_2007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2009 = 7'h2f == _myNewVec_113_T_3[6:0] ? myVec_47 : _GEN_2008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2010 = 7'h30 == _myNewVec_113_T_3[6:0] ? myVec_48 : _GEN_2009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2011 = 7'h31 == _myNewVec_113_T_3[6:0] ? myVec_49 : _GEN_2010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2012 = 7'h32 == _myNewVec_113_T_3[6:0] ? myVec_50 : _GEN_2011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2013 = 7'h33 == _myNewVec_113_T_3[6:0] ? myVec_51 : _GEN_2012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2014 = 7'h34 == _myNewVec_113_T_3[6:0] ? myVec_52 : _GEN_2013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2015 = 7'h35 == _myNewVec_113_T_3[6:0] ? myVec_53 : _GEN_2014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2016 = 7'h36 == _myNewVec_113_T_3[6:0] ? myVec_54 : _GEN_2015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2017 = 7'h37 == _myNewVec_113_T_3[6:0] ? myVec_55 : _GEN_2016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2018 = 7'h38 == _myNewVec_113_T_3[6:0] ? myVec_56 : _GEN_2017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2019 = 7'h39 == _myNewVec_113_T_3[6:0] ? myVec_57 : _GEN_2018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2020 = 7'h3a == _myNewVec_113_T_3[6:0] ? myVec_58 : _GEN_2019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2021 = 7'h3b == _myNewVec_113_T_3[6:0] ? myVec_59 : _GEN_2020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2022 = 7'h3c == _myNewVec_113_T_3[6:0] ? myVec_60 : _GEN_2021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2023 = 7'h3d == _myNewVec_113_T_3[6:0] ? myVec_61 : _GEN_2022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2024 = 7'h3e == _myNewVec_113_T_3[6:0] ? myVec_62 : _GEN_2023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2025 = 7'h3f == _myNewVec_113_T_3[6:0] ? myVec_63 : _GEN_2024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2026 = 7'h40 == _myNewVec_113_T_3[6:0] ? myVec_64 : _GEN_2025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2027 = 7'h41 == _myNewVec_113_T_3[6:0] ? myVec_65 : _GEN_2026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2028 = 7'h42 == _myNewVec_113_T_3[6:0] ? myVec_66 : _GEN_2027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2029 = 7'h43 == _myNewVec_113_T_3[6:0] ? myVec_67 : _GEN_2028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2030 = 7'h44 == _myNewVec_113_T_3[6:0] ? myVec_68 : _GEN_2029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2031 = 7'h45 == _myNewVec_113_T_3[6:0] ? myVec_69 : _GEN_2030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2032 = 7'h46 == _myNewVec_113_T_3[6:0] ? myVec_70 : _GEN_2031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2033 = 7'h47 == _myNewVec_113_T_3[6:0] ? myVec_71 : _GEN_2032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2034 = 7'h48 == _myNewVec_113_T_3[6:0] ? myVec_72 : _GEN_2033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2035 = 7'h49 == _myNewVec_113_T_3[6:0] ? myVec_73 : _GEN_2034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2036 = 7'h4a == _myNewVec_113_T_3[6:0] ? myVec_74 : _GEN_2035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2037 = 7'h4b == _myNewVec_113_T_3[6:0] ? myVec_75 : _GEN_2036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2038 = 7'h4c == _myNewVec_113_T_3[6:0] ? myVec_76 : _GEN_2037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2039 = 7'h4d == _myNewVec_113_T_3[6:0] ? myVec_77 : _GEN_2038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2040 = 7'h4e == _myNewVec_113_T_3[6:0] ? myVec_78 : _GEN_2039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2041 = 7'h4f == _myNewVec_113_T_3[6:0] ? myVec_79 : _GEN_2040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2042 = 7'h50 == _myNewVec_113_T_3[6:0] ? myVec_80 : _GEN_2041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2043 = 7'h51 == _myNewVec_113_T_3[6:0] ? myVec_81 : _GEN_2042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2044 = 7'h52 == _myNewVec_113_T_3[6:0] ? myVec_82 : _GEN_2043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2045 = 7'h53 == _myNewVec_113_T_3[6:0] ? myVec_83 : _GEN_2044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2046 = 7'h54 == _myNewVec_113_T_3[6:0] ? myVec_84 : _GEN_2045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2047 = 7'h55 == _myNewVec_113_T_3[6:0] ? myVec_85 : _GEN_2046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2048 = 7'h56 == _myNewVec_113_T_3[6:0] ? myVec_86 : _GEN_2047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2049 = 7'h57 == _myNewVec_113_T_3[6:0] ? myVec_87 : _GEN_2048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2050 = 7'h58 == _myNewVec_113_T_3[6:0] ? myVec_88 : _GEN_2049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2051 = 7'h59 == _myNewVec_113_T_3[6:0] ? myVec_89 : _GEN_2050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2052 = 7'h5a == _myNewVec_113_T_3[6:0] ? myVec_90 : _GEN_2051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2053 = 7'h5b == _myNewVec_113_T_3[6:0] ? myVec_91 : _GEN_2052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2054 = 7'h5c == _myNewVec_113_T_3[6:0] ? myVec_92 : _GEN_2053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2055 = 7'h5d == _myNewVec_113_T_3[6:0] ? myVec_93 : _GEN_2054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2056 = 7'h5e == _myNewVec_113_T_3[6:0] ? myVec_94 : _GEN_2055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2057 = 7'h5f == _myNewVec_113_T_3[6:0] ? myVec_95 : _GEN_2056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2058 = 7'h60 == _myNewVec_113_T_3[6:0] ? myVec_96 : _GEN_2057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2059 = 7'h61 == _myNewVec_113_T_3[6:0] ? myVec_97 : _GEN_2058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2060 = 7'h62 == _myNewVec_113_T_3[6:0] ? myVec_98 : _GEN_2059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2061 = 7'h63 == _myNewVec_113_T_3[6:0] ? myVec_99 : _GEN_2060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2062 = 7'h64 == _myNewVec_113_T_3[6:0] ? myVec_100 : _GEN_2061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2063 = 7'h65 == _myNewVec_113_T_3[6:0] ? myVec_101 : _GEN_2062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2064 = 7'h66 == _myNewVec_113_T_3[6:0] ? myVec_102 : _GEN_2063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2065 = 7'h67 == _myNewVec_113_T_3[6:0] ? myVec_103 : _GEN_2064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2066 = 7'h68 == _myNewVec_113_T_3[6:0] ? myVec_104 : _GEN_2065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2067 = 7'h69 == _myNewVec_113_T_3[6:0] ? myVec_105 : _GEN_2066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2068 = 7'h6a == _myNewVec_113_T_3[6:0] ? myVec_106 : _GEN_2067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2069 = 7'h6b == _myNewVec_113_T_3[6:0] ? myVec_107 : _GEN_2068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2070 = 7'h6c == _myNewVec_113_T_3[6:0] ? myVec_108 : _GEN_2069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2071 = 7'h6d == _myNewVec_113_T_3[6:0] ? myVec_109 : _GEN_2070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2072 = 7'h6e == _myNewVec_113_T_3[6:0] ? myVec_110 : _GEN_2071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2073 = 7'h6f == _myNewVec_113_T_3[6:0] ? myVec_111 : _GEN_2072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2074 = 7'h70 == _myNewVec_113_T_3[6:0] ? myVec_112 : _GEN_2073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2075 = 7'h71 == _myNewVec_113_T_3[6:0] ? myVec_113 : _GEN_2074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2076 = 7'h72 == _myNewVec_113_T_3[6:0] ? myVec_114 : _GEN_2075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2077 = 7'h73 == _myNewVec_113_T_3[6:0] ? myVec_115 : _GEN_2076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2078 = 7'h74 == _myNewVec_113_T_3[6:0] ? myVec_116 : _GEN_2077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2079 = 7'h75 == _myNewVec_113_T_3[6:0] ? myVec_117 : _GEN_2078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2080 = 7'h76 == _myNewVec_113_T_3[6:0] ? myVec_118 : _GEN_2079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2081 = 7'h77 == _myNewVec_113_T_3[6:0] ? myVec_119 : _GEN_2080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2082 = 7'h78 == _myNewVec_113_T_3[6:0] ? myVec_120 : _GEN_2081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2083 = 7'h79 == _myNewVec_113_T_3[6:0] ? myVec_121 : _GEN_2082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2084 = 7'h7a == _myNewVec_113_T_3[6:0] ? myVec_122 : _GEN_2083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2085 = 7'h7b == _myNewVec_113_T_3[6:0] ? myVec_123 : _GEN_2084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2086 = 7'h7c == _myNewVec_113_T_3[6:0] ? myVec_124 : _GEN_2085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2087 = 7'h7d == _myNewVec_113_T_3[6:0] ? myVec_125 : _GEN_2086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2088 = 7'h7e == _myNewVec_113_T_3[6:0] ? myVec_126 : _GEN_2087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_113 = 7'h7f == _myNewVec_113_T_3[6:0] ? myVec_127 : _GEN_2088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_112_T_3 = _myNewVec_127_T_1 + 16'hf; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2091 = 7'h1 == _myNewVec_112_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2092 = 7'h2 == _myNewVec_112_T_3[6:0] ? myVec_2 : _GEN_2091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2093 = 7'h3 == _myNewVec_112_T_3[6:0] ? myVec_3 : _GEN_2092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2094 = 7'h4 == _myNewVec_112_T_3[6:0] ? myVec_4 : _GEN_2093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2095 = 7'h5 == _myNewVec_112_T_3[6:0] ? myVec_5 : _GEN_2094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2096 = 7'h6 == _myNewVec_112_T_3[6:0] ? myVec_6 : _GEN_2095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2097 = 7'h7 == _myNewVec_112_T_3[6:0] ? myVec_7 : _GEN_2096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2098 = 7'h8 == _myNewVec_112_T_3[6:0] ? myVec_8 : _GEN_2097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2099 = 7'h9 == _myNewVec_112_T_3[6:0] ? myVec_9 : _GEN_2098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2100 = 7'ha == _myNewVec_112_T_3[6:0] ? myVec_10 : _GEN_2099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2101 = 7'hb == _myNewVec_112_T_3[6:0] ? myVec_11 : _GEN_2100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2102 = 7'hc == _myNewVec_112_T_3[6:0] ? myVec_12 : _GEN_2101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2103 = 7'hd == _myNewVec_112_T_3[6:0] ? myVec_13 : _GEN_2102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2104 = 7'he == _myNewVec_112_T_3[6:0] ? myVec_14 : _GEN_2103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2105 = 7'hf == _myNewVec_112_T_3[6:0] ? myVec_15 : _GEN_2104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2106 = 7'h10 == _myNewVec_112_T_3[6:0] ? myVec_16 : _GEN_2105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2107 = 7'h11 == _myNewVec_112_T_3[6:0] ? myVec_17 : _GEN_2106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2108 = 7'h12 == _myNewVec_112_T_3[6:0] ? myVec_18 : _GEN_2107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2109 = 7'h13 == _myNewVec_112_T_3[6:0] ? myVec_19 : _GEN_2108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2110 = 7'h14 == _myNewVec_112_T_3[6:0] ? myVec_20 : _GEN_2109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2111 = 7'h15 == _myNewVec_112_T_3[6:0] ? myVec_21 : _GEN_2110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2112 = 7'h16 == _myNewVec_112_T_3[6:0] ? myVec_22 : _GEN_2111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2113 = 7'h17 == _myNewVec_112_T_3[6:0] ? myVec_23 : _GEN_2112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2114 = 7'h18 == _myNewVec_112_T_3[6:0] ? myVec_24 : _GEN_2113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2115 = 7'h19 == _myNewVec_112_T_3[6:0] ? myVec_25 : _GEN_2114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2116 = 7'h1a == _myNewVec_112_T_3[6:0] ? myVec_26 : _GEN_2115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2117 = 7'h1b == _myNewVec_112_T_3[6:0] ? myVec_27 : _GEN_2116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2118 = 7'h1c == _myNewVec_112_T_3[6:0] ? myVec_28 : _GEN_2117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2119 = 7'h1d == _myNewVec_112_T_3[6:0] ? myVec_29 : _GEN_2118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2120 = 7'h1e == _myNewVec_112_T_3[6:0] ? myVec_30 : _GEN_2119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2121 = 7'h1f == _myNewVec_112_T_3[6:0] ? myVec_31 : _GEN_2120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2122 = 7'h20 == _myNewVec_112_T_3[6:0] ? myVec_32 : _GEN_2121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2123 = 7'h21 == _myNewVec_112_T_3[6:0] ? myVec_33 : _GEN_2122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2124 = 7'h22 == _myNewVec_112_T_3[6:0] ? myVec_34 : _GEN_2123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2125 = 7'h23 == _myNewVec_112_T_3[6:0] ? myVec_35 : _GEN_2124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2126 = 7'h24 == _myNewVec_112_T_3[6:0] ? myVec_36 : _GEN_2125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2127 = 7'h25 == _myNewVec_112_T_3[6:0] ? myVec_37 : _GEN_2126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2128 = 7'h26 == _myNewVec_112_T_3[6:0] ? myVec_38 : _GEN_2127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2129 = 7'h27 == _myNewVec_112_T_3[6:0] ? myVec_39 : _GEN_2128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2130 = 7'h28 == _myNewVec_112_T_3[6:0] ? myVec_40 : _GEN_2129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2131 = 7'h29 == _myNewVec_112_T_3[6:0] ? myVec_41 : _GEN_2130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2132 = 7'h2a == _myNewVec_112_T_3[6:0] ? myVec_42 : _GEN_2131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2133 = 7'h2b == _myNewVec_112_T_3[6:0] ? myVec_43 : _GEN_2132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2134 = 7'h2c == _myNewVec_112_T_3[6:0] ? myVec_44 : _GEN_2133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2135 = 7'h2d == _myNewVec_112_T_3[6:0] ? myVec_45 : _GEN_2134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2136 = 7'h2e == _myNewVec_112_T_3[6:0] ? myVec_46 : _GEN_2135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2137 = 7'h2f == _myNewVec_112_T_3[6:0] ? myVec_47 : _GEN_2136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2138 = 7'h30 == _myNewVec_112_T_3[6:0] ? myVec_48 : _GEN_2137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2139 = 7'h31 == _myNewVec_112_T_3[6:0] ? myVec_49 : _GEN_2138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2140 = 7'h32 == _myNewVec_112_T_3[6:0] ? myVec_50 : _GEN_2139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2141 = 7'h33 == _myNewVec_112_T_3[6:0] ? myVec_51 : _GEN_2140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2142 = 7'h34 == _myNewVec_112_T_3[6:0] ? myVec_52 : _GEN_2141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2143 = 7'h35 == _myNewVec_112_T_3[6:0] ? myVec_53 : _GEN_2142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2144 = 7'h36 == _myNewVec_112_T_3[6:0] ? myVec_54 : _GEN_2143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2145 = 7'h37 == _myNewVec_112_T_3[6:0] ? myVec_55 : _GEN_2144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2146 = 7'h38 == _myNewVec_112_T_3[6:0] ? myVec_56 : _GEN_2145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2147 = 7'h39 == _myNewVec_112_T_3[6:0] ? myVec_57 : _GEN_2146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2148 = 7'h3a == _myNewVec_112_T_3[6:0] ? myVec_58 : _GEN_2147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2149 = 7'h3b == _myNewVec_112_T_3[6:0] ? myVec_59 : _GEN_2148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2150 = 7'h3c == _myNewVec_112_T_3[6:0] ? myVec_60 : _GEN_2149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2151 = 7'h3d == _myNewVec_112_T_3[6:0] ? myVec_61 : _GEN_2150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2152 = 7'h3e == _myNewVec_112_T_3[6:0] ? myVec_62 : _GEN_2151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2153 = 7'h3f == _myNewVec_112_T_3[6:0] ? myVec_63 : _GEN_2152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2154 = 7'h40 == _myNewVec_112_T_3[6:0] ? myVec_64 : _GEN_2153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2155 = 7'h41 == _myNewVec_112_T_3[6:0] ? myVec_65 : _GEN_2154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2156 = 7'h42 == _myNewVec_112_T_3[6:0] ? myVec_66 : _GEN_2155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2157 = 7'h43 == _myNewVec_112_T_3[6:0] ? myVec_67 : _GEN_2156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2158 = 7'h44 == _myNewVec_112_T_3[6:0] ? myVec_68 : _GEN_2157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2159 = 7'h45 == _myNewVec_112_T_3[6:0] ? myVec_69 : _GEN_2158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2160 = 7'h46 == _myNewVec_112_T_3[6:0] ? myVec_70 : _GEN_2159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2161 = 7'h47 == _myNewVec_112_T_3[6:0] ? myVec_71 : _GEN_2160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2162 = 7'h48 == _myNewVec_112_T_3[6:0] ? myVec_72 : _GEN_2161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2163 = 7'h49 == _myNewVec_112_T_3[6:0] ? myVec_73 : _GEN_2162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2164 = 7'h4a == _myNewVec_112_T_3[6:0] ? myVec_74 : _GEN_2163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2165 = 7'h4b == _myNewVec_112_T_3[6:0] ? myVec_75 : _GEN_2164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2166 = 7'h4c == _myNewVec_112_T_3[6:0] ? myVec_76 : _GEN_2165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2167 = 7'h4d == _myNewVec_112_T_3[6:0] ? myVec_77 : _GEN_2166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2168 = 7'h4e == _myNewVec_112_T_3[6:0] ? myVec_78 : _GEN_2167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2169 = 7'h4f == _myNewVec_112_T_3[6:0] ? myVec_79 : _GEN_2168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2170 = 7'h50 == _myNewVec_112_T_3[6:0] ? myVec_80 : _GEN_2169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2171 = 7'h51 == _myNewVec_112_T_3[6:0] ? myVec_81 : _GEN_2170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2172 = 7'h52 == _myNewVec_112_T_3[6:0] ? myVec_82 : _GEN_2171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2173 = 7'h53 == _myNewVec_112_T_3[6:0] ? myVec_83 : _GEN_2172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2174 = 7'h54 == _myNewVec_112_T_3[6:0] ? myVec_84 : _GEN_2173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2175 = 7'h55 == _myNewVec_112_T_3[6:0] ? myVec_85 : _GEN_2174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2176 = 7'h56 == _myNewVec_112_T_3[6:0] ? myVec_86 : _GEN_2175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2177 = 7'h57 == _myNewVec_112_T_3[6:0] ? myVec_87 : _GEN_2176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2178 = 7'h58 == _myNewVec_112_T_3[6:0] ? myVec_88 : _GEN_2177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2179 = 7'h59 == _myNewVec_112_T_3[6:0] ? myVec_89 : _GEN_2178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2180 = 7'h5a == _myNewVec_112_T_3[6:0] ? myVec_90 : _GEN_2179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2181 = 7'h5b == _myNewVec_112_T_3[6:0] ? myVec_91 : _GEN_2180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2182 = 7'h5c == _myNewVec_112_T_3[6:0] ? myVec_92 : _GEN_2181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2183 = 7'h5d == _myNewVec_112_T_3[6:0] ? myVec_93 : _GEN_2182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2184 = 7'h5e == _myNewVec_112_T_3[6:0] ? myVec_94 : _GEN_2183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2185 = 7'h5f == _myNewVec_112_T_3[6:0] ? myVec_95 : _GEN_2184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2186 = 7'h60 == _myNewVec_112_T_3[6:0] ? myVec_96 : _GEN_2185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2187 = 7'h61 == _myNewVec_112_T_3[6:0] ? myVec_97 : _GEN_2186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2188 = 7'h62 == _myNewVec_112_T_3[6:0] ? myVec_98 : _GEN_2187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2189 = 7'h63 == _myNewVec_112_T_3[6:0] ? myVec_99 : _GEN_2188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2190 = 7'h64 == _myNewVec_112_T_3[6:0] ? myVec_100 : _GEN_2189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2191 = 7'h65 == _myNewVec_112_T_3[6:0] ? myVec_101 : _GEN_2190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2192 = 7'h66 == _myNewVec_112_T_3[6:0] ? myVec_102 : _GEN_2191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2193 = 7'h67 == _myNewVec_112_T_3[6:0] ? myVec_103 : _GEN_2192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2194 = 7'h68 == _myNewVec_112_T_3[6:0] ? myVec_104 : _GEN_2193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2195 = 7'h69 == _myNewVec_112_T_3[6:0] ? myVec_105 : _GEN_2194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2196 = 7'h6a == _myNewVec_112_T_3[6:0] ? myVec_106 : _GEN_2195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2197 = 7'h6b == _myNewVec_112_T_3[6:0] ? myVec_107 : _GEN_2196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2198 = 7'h6c == _myNewVec_112_T_3[6:0] ? myVec_108 : _GEN_2197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2199 = 7'h6d == _myNewVec_112_T_3[6:0] ? myVec_109 : _GEN_2198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2200 = 7'h6e == _myNewVec_112_T_3[6:0] ? myVec_110 : _GEN_2199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2201 = 7'h6f == _myNewVec_112_T_3[6:0] ? myVec_111 : _GEN_2200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2202 = 7'h70 == _myNewVec_112_T_3[6:0] ? myVec_112 : _GEN_2201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2203 = 7'h71 == _myNewVec_112_T_3[6:0] ? myVec_113 : _GEN_2202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2204 = 7'h72 == _myNewVec_112_T_3[6:0] ? myVec_114 : _GEN_2203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2205 = 7'h73 == _myNewVec_112_T_3[6:0] ? myVec_115 : _GEN_2204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2206 = 7'h74 == _myNewVec_112_T_3[6:0] ? myVec_116 : _GEN_2205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2207 = 7'h75 == _myNewVec_112_T_3[6:0] ? myVec_117 : _GEN_2206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2208 = 7'h76 == _myNewVec_112_T_3[6:0] ? myVec_118 : _GEN_2207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2209 = 7'h77 == _myNewVec_112_T_3[6:0] ? myVec_119 : _GEN_2208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2210 = 7'h78 == _myNewVec_112_T_3[6:0] ? myVec_120 : _GEN_2209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2211 = 7'h79 == _myNewVec_112_T_3[6:0] ? myVec_121 : _GEN_2210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2212 = 7'h7a == _myNewVec_112_T_3[6:0] ? myVec_122 : _GEN_2211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2213 = 7'h7b == _myNewVec_112_T_3[6:0] ? myVec_123 : _GEN_2212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2214 = 7'h7c == _myNewVec_112_T_3[6:0] ? myVec_124 : _GEN_2213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2215 = 7'h7d == _myNewVec_112_T_3[6:0] ? myVec_125 : _GEN_2214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2216 = 7'h7e == _myNewVec_112_T_3[6:0] ? myVec_126 : _GEN_2215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_112 = 7'h7f == _myNewVec_112_T_3[6:0] ? myVec_127 : _GEN_2216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [255:0] myNewWire_hi_hi_hi_lo = {myNewVec_119,myNewVec_118,myNewVec_117,myNewVec_116,myNewVec_115,myNewVec_114,
    myNewVec_113,myNewVec_112}; // @[hh_datapath_chisel.scala 238:27]
  wire [15:0] _myNewVec_111_T_3 = _myNewVec_127_T_1 + 16'h10; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2219 = 7'h1 == _myNewVec_111_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2220 = 7'h2 == _myNewVec_111_T_3[6:0] ? myVec_2 : _GEN_2219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2221 = 7'h3 == _myNewVec_111_T_3[6:0] ? myVec_3 : _GEN_2220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2222 = 7'h4 == _myNewVec_111_T_3[6:0] ? myVec_4 : _GEN_2221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2223 = 7'h5 == _myNewVec_111_T_3[6:0] ? myVec_5 : _GEN_2222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2224 = 7'h6 == _myNewVec_111_T_3[6:0] ? myVec_6 : _GEN_2223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2225 = 7'h7 == _myNewVec_111_T_3[6:0] ? myVec_7 : _GEN_2224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2226 = 7'h8 == _myNewVec_111_T_3[6:0] ? myVec_8 : _GEN_2225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2227 = 7'h9 == _myNewVec_111_T_3[6:0] ? myVec_9 : _GEN_2226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2228 = 7'ha == _myNewVec_111_T_3[6:0] ? myVec_10 : _GEN_2227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2229 = 7'hb == _myNewVec_111_T_3[6:0] ? myVec_11 : _GEN_2228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2230 = 7'hc == _myNewVec_111_T_3[6:0] ? myVec_12 : _GEN_2229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2231 = 7'hd == _myNewVec_111_T_3[6:0] ? myVec_13 : _GEN_2230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2232 = 7'he == _myNewVec_111_T_3[6:0] ? myVec_14 : _GEN_2231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2233 = 7'hf == _myNewVec_111_T_3[6:0] ? myVec_15 : _GEN_2232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2234 = 7'h10 == _myNewVec_111_T_3[6:0] ? myVec_16 : _GEN_2233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2235 = 7'h11 == _myNewVec_111_T_3[6:0] ? myVec_17 : _GEN_2234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2236 = 7'h12 == _myNewVec_111_T_3[6:0] ? myVec_18 : _GEN_2235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2237 = 7'h13 == _myNewVec_111_T_3[6:0] ? myVec_19 : _GEN_2236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2238 = 7'h14 == _myNewVec_111_T_3[6:0] ? myVec_20 : _GEN_2237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2239 = 7'h15 == _myNewVec_111_T_3[6:0] ? myVec_21 : _GEN_2238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2240 = 7'h16 == _myNewVec_111_T_3[6:0] ? myVec_22 : _GEN_2239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2241 = 7'h17 == _myNewVec_111_T_3[6:0] ? myVec_23 : _GEN_2240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2242 = 7'h18 == _myNewVec_111_T_3[6:0] ? myVec_24 : _GEN_2241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2243 = 7'h19 == _myNewVec_111_T_3[6:0] ? myVec_25 : _GEN_2242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2244 = 7'h1a == _myNewVec_111_T_3[6:0] ? myVec_26 : _GEN_2243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2245 = 7'h1b == _myNewVec_111_T_3[6:0] ? myVec_27 : _GEN_2244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2246 = 7'h1c == _myNewVec_111_T_3[6:0] ? myVec_28 : _GEN_2245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2247 = 7'h1d == _myNewVec_111_T_3[6:0] ? myVec_29 : _GEN_2246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2248 = 7'h1e == _myNewVec_111_T_3[6:0] ? myVec_30 : _GEN_2247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2249 = 7'h1f == _myNewVec_111_T_3[6:0] ? myVec_31 : _GEN_2248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2250 = 7'h20 == _myNewVec_111_T_3[6:0] ? myVec_32 : _GEN_2249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2251 = 7'h21 == _myNewVec_111_T_3[6:0] ? myVec_33 : _GEN_2250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2252 = 7'h22 == _myNewVec_111_T_3[6:0] ? myVec_34 : _GEN_2251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2253 = 7'h23 == _myNewVec_111_T_3[6:0] ? myVec_35 : _GEN_2252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2254 = 7'h24 == _myNewVec_111_T_3[6:0] ? myVec_36 : _GEN_2253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2255 = 7'h25 == _myNewVec_111_T_3[6:0] ? myVec_37 : _GEN_2254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2256 = 7'h26 == _myNewVec_111_T_3[6:0] ? myVec_38 : _GEN_2255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2257 = 7'h27 == _myNewVec_111_T_3[6:0] ? myVec_39 : _GEN_2256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2258 = 7'h28 == _myNewVec_111_T_3[6:0] ? myVec_40 : _GEN_2257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2259 = 7'h29 == _myNewVec_111_T_3[6:0] ? myVec_41 : _GEN_2258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2260 = 7'h2a == _myNewVec_111_T_3[6:0] ? myVec_42 : _GEN_2259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2261 = 7'h2b == _myNewVec_111_T_3[6:0] ? myVec_43 : _GEN_2260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2262 = 7'h2c == _myNewVec_111_T_3[6:0] ? myVec_44 : _GEN_2261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2263 = 7'h2d == _myNewVec_111_T_3[6:0] ? myVec_45 : _GEN_2262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2264 = 7'h2e == _myNewVec_111_T_3[6:0] ? myVec_46 : _GEN_2263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2265 = 7'h2f == _myNewVec_111_T_3[6:0] ? myVec_47 : _GEN_2264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2266 = 7'h30 == _myNewVec_111_T_3[6:0] ? myVec_48 : _GEN_2265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2267 = 7'h31 == _myNewVec_111_T_3[6:0] ? myVec_49 : _GEN_2266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2268 = 7'h32 == _myNewVec_111_T_3[6:0] ? myVec_50 : _GEN_2267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2269 = 7'h33 == _myNewVec_111_T_3[6:0] ? myVec_51 : _GEN_2268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2270 = 7'h34 == _myNewVec_111_T_3[6:0] ? myVec_52 : _GEN_2269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2271 = 7'h35 == _myNewVec_111_T_3[6:0] ? myVec_53 : _GEN_2270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2272 = 7'h36 == _myNewVec_111_T_3[6:0] ? myVec_54 : _GEN_2271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2273 = 7'h37 == _myNewVec_111_T_3[6:0] ? myVec_55 : _GEN_2272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2274 = 7'h38 == _myNewVec_111_T_3[6:0] ? myVec_56 : _GEN_2273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2275 = 7'h39 == _myNewVec_111_T_3[6:0] ? myVec_57 : _GEN_2274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2276 = 7'h3a == _myNewVec_111_T_3[6:0] ? myVec_58 : _GEN_2275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2277 = 7'h3b == _myNewVec_111_T_3[6:0] ? myVec_59 : _GEN_2276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2278 = 7'h3c == _myNewVec_111_T_3[6:0] ? myVec_60 : _GEN_2277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2279 = 7'h3d == _myNewVec_111_T_3[6:0] ? myVec_61 : _GEN_2278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2280 = 7'h3e == _myNewVec_111_T_3[6:0] ? myVec_62 : _GEN_2279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2281 = 7'h3f == _myNewVec_111_T_3[6:0] ? myVec_63 : _GEN_2280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2282 = 7'h40 == _myNewVec_111_T_3[6:0] ? myVec_64 : _GEN_2281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2283 = 7'h41 == _myNewVec_111_T_3[6:0] ? myVec_65 : _GEN_2282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2284 = 7'h42 == _myNewVec_111_T_3[6:0] ? myVec_66 : _GEN_2283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2285 = 7'h43 == _myNewVec_111_T_3[6:0] ? myVec_67 : _GEN_2284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2286 = 7'h44 == _myNewVec_111_T_3[6:0] ? myVec_68 : _GEN_2285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2287 = 7'h45 == _myNewVec_111_T_3[6:0] ? myVec_69 : _GEN_2286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2288 = 7'h46 == _myNewVec_111_T_3[6:0] ? myVec_70 : _GEN_2287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2289 = 7'h47 == _myNewVec_111_T_3[6:0] ? myVec_71 : _GEN_2288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2290 = 7'h48 == _myNewVec_111_T_3[6:0] ? myVec_72 : _GEN_2289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2291 = 7'h49 == _myNewVec_111_T_3[6:0] ? myVec_73 : _GEN_2290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2292 = 7'h4a == _myNewVec_111_T_3[6:0] ? myVec_74 : _GEN_2291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2293 = 7'h4b == _myNewVec_111_T_3[6:0] ? myVec_75 : _GEN_2292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2294 = 7'h4c == _myNewVec_111_T_3[6:0] ? myVec_76 : _GEN_2293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2295 = 7'h4d == _myNewVec_111_T_3[6:0] ? myVec_77 : _GEN_2294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2296 = 7'h4e == _myNewVec_111_T_3[6:0] ? myVec_78 : _GEN_2295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2297 = 7'h4f == _myNewVec_111_T_3[6:0] ? myVec_79 : _GEN_2296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2298 = 7'h50 == _myNewVec_111_T_3[6:0] ? myVec_80 : _GEN_2297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2299 = 7'h51 == _myNewVec_111_T_3[6:0] ? myVec_81 : _GEN_2298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2300 = 7'h52 == _myNewVec_111_T_3[6:0] ? myVec_82 : _GEN_2299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2301 = 7'h53 == _myNewVec_111_T_3[6:0] ? myVec_83 : _GEN_2300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2302 = 7'h54 == _myNewVec_111_T_3[6:0] ? myVec_84 : _GEN_2301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2303 = 7'h55 == _myNewVec_111_T_3[6:0] ? myVec_85 : _GEN_2302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2304 = 7'h56 == _myNewVec_111_T_3[6:0] ? myVec_86 : _GEN_2303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2305 = 7'h57 == _myNewVec_111_T_3[6:0] ? myVec_87 : _GEN_2304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2306 = 7'h58 == _myNewVec_111_T_3[6:0] ? myVec_88 : _GEN_2305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2307 = 7'h59 == _myNewVec_111_T_3[6:0] ? myVec_89 : _GEN_2306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2308 = 7'h5a == _myNewVec_111_T_3[6:0] ? myVec_90 : _GEN_2307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2309 = 7'h5b == _myNewVec_111_T_3[6:0] ? myVec_91 : _GEN_2308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2310 = 7'h5c == _myNewVec_111_T_3[6:0] ? myVec_92 : _GEN_2309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2311 = 7'h5d == _myNewVec_111_T_3[6:0] ? myVec_93 : _GEN_2310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2312 = 7'h5e == _myNewVec_111_T_3[6:0] ? myVec_94 : _GEN_2311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2313 = 7'h5f == _myNewVec_111_T_3[6:0] ? myVec_95 : _GEN_2312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2314 = 7'h60 == _myNewVec_111_T_3[6:0] ? myVec_96 : _GEN_2313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2315 = 7'h61 == _myNewVec_111_T_3[6:0] ? myVec_97 : _GEN_2314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2316 = 7'h62 == _myNewVec_111_T_3[6:0] ? myVec_98 : _GEN_2315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2317 = 7'h63 == _myNewVec_111_T_3[6:0] ? myVec_99 : _GEN_2316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2318 = 7'h64 == _myNewVec_111_T_3[6:0] ? myVec_100 : _GEN_2317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2319 = 7'h65 == _myNewVec_111_T_3[6:0] ? myVec_101 : _GEN_2318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2320 = 7'h66 == _myNewVec_111_T_3[6:0] ? myVec_102 : _GEN_2319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2321 = 7'h67 == _myNewVec_111_T_3[6:0] ? myVec_103 : _GEN_2320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2322 = 7'h68 == _myNewVec_111_T_3[6:0] ? myVec_104 : _GEN_2321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2323 = 7'h69 == _myNewVec_111_T_3[6:0] ? myVec_105 : _GEN_2322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2324 = 7'h6a == _myNewVec_111_T_3[6:0] ? myVec_106 : _GEN_2323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2325 = 7'h6b == _myNewVec_111_T_3[6:0] ? myVec_107 : _GEN_2324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2326 = 7'h6c == _myNewVec_111_T_3[6:0] ? myVec_108 : _GEN_2325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2327 = 7'h6d == _myNewVec_111_T_3[6:0] ? myVec_109 : _GEN_2326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2328 = 7'h6e == _myNewVec_111_T_3[6:0] ? myVec_110 : _GEN_2327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2329 = 7'h6f == _myNewVec_111_T_3[6:0] ? myVec_111 : _GEN_2328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2330 = 7'h70 == _myNewVec_111_T_3[6:0] ? myVec_112 : _GEN_2329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2331 = 7'h71 == _myNewVec_111_T_3[6:0] ? myVec_113 : _GEN_2330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2332 = 7'h72 == _myNewVec_111_T_3[6:0] ? myVec_114 : _GEN_2331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2333 = 7'h73 == _myNewVec_111_T_3[6:0] ? myVec_115 : _GEN_2332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2334 = 7'h74 == _myNewVec_111_T_3[6:0] ? myVec_116 : _GEN_2333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2335 = 7'h75 == _myNewVec_111_T_3[6:0] ? myVec_117 : _GEN_2334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2336 = 7'h76 == _myNewVec_111_T_3[6:0] ? myVec_118 : _GEN_2335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2337 = 7'h77 == _myNewVec_111_T_3[6:0] ? myVec_119 : _GEN_2336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2338 = 7'h78 == _myNewVec_111_T_3[6:0] ? myVec_120 : _GEN_2337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2339 = 7'h79 == _myNewVec_111_T_3[6:0] ? myVec_121 : _GEN_2338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2340 = 7'h7a == _myNewVec_111_T_3[6:0] ? myVec_122 : _GEN_2339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2341 = 7'h7b == _myNewVec_111_T_3[6:0] ? myVec_123 : _GEN_2340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2342 = 7'h7c == _myNewVec_111_T_3[6:0] ? myVec_124 : _GEN_2341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2343 = 7'h7d == _myNewVec_111_T_3[6:0] ? myVec_125 : _GEN_2342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2344 = 7'h7e == _myNewVec_111_T_3[6:0] ? myVec_126 : _GEN_2343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_111 = 7'h7f == _myNewVec_111_T_3[6:0] ? myVec_127 : _GEN_2344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_110_T_3 = _myNewVec_127_T_1 + 16'h11; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2347 = 7'h1 == _myNewVec_110_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2348 = 7'h2 == _myNewVec_110_T_3[6:0] ? myVec_2 : _GEN_2347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2349 = 7'h3 == _myNewVec_110_T_3[6:0] ? myVec_3 : _GEN_2348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2350 = 7'h4 == _myNewVec_110_T_3[6:0] ? myVec_4 : _GEN_2349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2351 = 7'h5 == _myNewVec_110_T_3[6:0] ? myVec_5 : _GEN_2350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2352 = 7'h6 == _myNewVec_110_T_3[6:0] ? myVec_6 : _GEN_2351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2353 = 7'h7 == _myNewVec_110_T_3[6:0] ? myVec_7 : _GEN_2352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2354 = 7'h8 == _myNewVec_110_T_3[6:0] ? myVec_8 : _GEN_2353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2355 = 7'h9 == _myNewVec_110_T_3[6:0] ? myVec_9 : _GEN_2354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2356 = 7'ha == _myNewVec_110_T_3[6:0] ? myVec_10 : _GEN_2355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2357 = 7'hb == _myNewVec_110_T_3[6:0] ? myVec_11 : _GEN_2356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2358 = 7'hc == _myNewVec_110_T_3[6:0] ? myVec_12 : _GEN_2357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2359 = 7'hd == _myNewVec_110_T_3[6:0] ? myVec_13 : _GEN_2358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2360 = 7'he == _myNewVec_110_T_3[6:0] ? myVec_14 : _GEN_2359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2361 = 7'hf == _myNewVec_110_T_3[6:0] ? myVec_15 : _GEN_2360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2362 = 7'h10 == _myNewVec_110_T_3[6:0] ? myVec_16 : _GEN_2361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2363 = 7'h11 == _myNewVec_110_T_3[6:0] ? myVec_17 : _GEN_2362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2364 = 7'h12 == _myNewVec_110_T_3[6:0] ? myVec_18 : _GEN_2363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2365 = 7'h13 == _myNewVec_110_T_3[6:0] ? myVec_19 : _GEN_2364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2366 = 7'h14 == _myNewVec_110_T_3[6:0] ? myVec_20 : _GEN_2365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2367 = 7'h15 == _myNewVec_110_T_3[6:0] ? myVec_21 : _GEN_2366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2368 = 7'h16 == _myNewVec_110_T_3[6:0] ? myVec_22 : _GEN_2367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2369 = 7'h17 == _myNewVec_110_T_3[6:0] ? myVec_23 : _GEN_2368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2370 = 7'h18 == _myNewVec_110_T_3[6:0] ? myVec_24 : _GEN_2369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2371 = 7'h19 == _myNewVec_110_T_3[6:0] ? myVec_25 : _GEN_2370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2372 = 7'h1a == _myNewVec_110_T_3[6:0] ? myVec_26 : _GEN_2371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2373 = 7'h1b == _myNewVec_110_T_3[6:0] ? myVec_27 : _GEN_2372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2374 = 7'h1c == _myNewVec_110_T_3[6:0] ? myVec_28 : _GEN_2373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2375 = 7'h1d == _myNewVec_110_T_3[6:0] ? myVec_29 : _GEN_2374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2376 = 7'h1e == _myNewVec_110_T_3[6:0] ? myVec_30 : _GEN_2375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2377 = 7'h1f == _myNewVec_110_T_3[6:0] ? myVec_31 : _GEN_2376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2378 = 7'h20 == _myNewVec_110_T_3[6:0] ? myVec_32 : _GEN_2377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2379 = 7'h21 == _myNewVec_110_T_3[6:0] ? myVec_33 : _GEN_2378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2380 = 7'h22 == _myNewVec_110_T_3[6:0] ? myVec_34 : _GEN_2379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2381 = 7'h23 == _myNewVec_110_T_3[6:0] ? myVec_35 : _GEN_2380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2382 = 7'h24 == _myNewVec_110_T_3[6:0] ? myVec_36 : _GEN_2381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2383 = 7'h25 == _myNewVec_110_T_3[6:0] ? myVec_37 : _GEN_2382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2384 = 7'h26 == _myNewVec_110_T_3[6:0] ? myVec_38 : _GEN_2383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2385 = 7'h27 == _myNewVec_110_T_3[6:0] ? myVec_39 : _GEN_2384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2386 = 7'h28 == _myNewVec_110_T_3[6:0] ? myVec_40 : _GEN_2385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2387 = 7'h29 == _myNewVec_110_T_3[6:0] ? myVec_41 : _GEN_2386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2388 = 7'h2a == _myNewVec_110_T_3[6:0] ? myVec_42 : _GEN_2387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2389 = 7'h2b == _myNewVec_110_T_3[6:0] ? myVec_43 : _GEN_2388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2390 = 7'h2c == _myNewVec_110_T_3[6:0] ? myVec_44 : _GEN_2389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2391 = 7'h2d == _myNewVec_110_T_3[6:0] ? myVec_45 : _GEN_2390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2392 = 7'h2e == _myNewVec_110_T_3[6:0] ? myVec_46 : _GEN_2391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2393 = 7'h2f == _myNewVec_110_T_3[6:0] ? myVec_47 : _GEN_2392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2394 = 7'h30 == _myNewVec_110_T_3[6:0] ? myVec_48 : _GEN_2393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2395 = 7'h31 == _myNewVec_110_T_3[6:0] ? myVec_49 : _GEN_2394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2396 = 7'h32 == _myNewVec_110_T_3[6:0] ? myVec_50 : _GEN_2395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2397 = 7'h33 == _myNewVec_110_T_3[6:0] ? myVec_51 : _GEN_2396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2398 = 7'h34 == _myNewVec_110_T_3[6:0] ? myVec_52 : _GEN_2397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2399 = 7'h35 == _myNewVec_110_T_3[6:0] ? myVec_53 : _GEN_2398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2400 = 7'h36 == _myNewVec_110_T_3[6:0] ? myVec_54 : _GEN_2399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2401 = 7'h37 == _myNewVec_110_T_3[6:0] ? myVec_55 : _GEN_2400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2402 = 7'h38 == _myNewVec_110_T_3[6:0] ? myVec_56 : _GEN_2401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2403 = 7'h39 == _myNewVec_110_T_3[6:0] ? myVec_57 : _GEN_2402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2404 = 7'h3a == _myNewVec_110_T_3[6:0] ? myVec_58 : _GEN_2403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2405 = 7'h3b == _myNewVec_110_T_3[6:0] ? myVec_59 : _GEN_2404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2406 = 7'h3c == _myNewVec_110_T_3[6:0] ? myVec_60 : _GEN_2405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2407 = 7'h3d == _myNewVec_110_T_3[6:0] ? myVec_61 : _GEN_2406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2408 = 7'h3e == _myNewVec_110_T_3[6:0] ? myVec_62 : _GEN_2407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2409 = 7'h3f == _myNewVec_110_T_3[6:0] ? myVec_63 : _GEN_2408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2410 = 7'h40 == _myNewVec_110_T_3[6:0] ? myVec_64 : _GEN_2409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2411 = 7'h41 == _myNewVec_110_T_3[6:0] ? myVec_65 : _GEN_2410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2412 = 7'h42 == _myNewVec_110_T_3[6:0] ? myVec_66 : _GEN_2411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2413 = 7'h43 == _myNewVec_110_T_3[6:0] ? myVec_67 : _GEN_2412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2414 = 7'h44 == _myNewVec_110_T_3[6:0] ? myVec_68 : _GEN_2413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2415 = 7'h45 == _myNewVec_110_T_3[6:0] ? myVec_69 : _GEN_2414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2416 = 7'h46 == _myNewVec_110_T_3[6:0] ? myVec_70 : _GEN_2415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2417 = 7'h47 == _myNewVec_110_T_3[6:0] ? myVec_71 : _GEN_2416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2418 = 7'h48 == _myNewVec_110_T_3[6:0] ? myVec_72 : _GEN_2417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2419 = 7'h49 == _myNewVec_110_T_3[6:0] ? myVec_73 : _GEN_2418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2420 = 7'h4a == _myNewVec_110_T_3[6:0] ? myVec_74 : _GEN_2419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2421 = 7'h4b == _myNewVec_110_T_3[6:0] ? myVec_75 : _GEN_2420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2422 = 7'h4c == _myNewVec_110_T_3[6:0] ? myVec_76 : _GEN_2421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2423 = 7'h4d == _myNewVec_110_T_3[6:0] ? myVec_77 : _GEN_2422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2424 = 7'h4e == _myNewVec_110_T_3[6:0] ? myVec_78 : _GEN_2423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2425 = 7'h4f == _myNewVec_110_T_3[6:0] ? myVec_79 : _GEN_2424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2426 = 7'h50 == _myNewVec_110_T_3[6:0] ? myVec_80 : _GEN_2425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2427 = 7'h51 == _myNewVec_110_T_3[6:0] ? myVec_81 : _GEN_2426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2428 = 7'h52 == _myNewVec_110_T_3[6:0] ? myVec_82 : _GEN_2427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2429 = 7'h53 == _myNewVec_110_T_3[6:0] ? myVec_83 : _GEN_2428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2430 = 7'h54 == _myNewVec_110_T_3[6:0] ? myVec_84 : _GEN_2429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2431 = 7'h55 == _myNewVec_110_T_3[6:0] ? myVec_85 : _GEN_2430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2432 = 7'h56 == _myNewVec_110_T_3[6:0] ? myVec_86 : _GEN_2431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2433 = 7'h57 == _myNewVec_110_T_3[6:0] ? myVec_87 : _GEN_2432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2434 = 7'h58 == _myNewVec_110_T_3[6:0] ? myVec_88 : _GEN_2433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2435 = 7'h59 == _myNewVec_110_T_3[6:0] ? myVec_89 : _GEN_2434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2436 = 7'h5a == _myNewVec_110_T_3[6:0] ? myVec_90 : _GEN_2435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2437 = 7'h5b == _myNewVec_110_T_3[6:0] ? myVec_91 : _GEN_2436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2438 = 7'h5c == _myNewVec_110_T_3[6:0] ? myVec_92 : _GEN_2437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2439 = 7'h5d == _myNewVec_110_T_3[6:0] ? myVec_93 : _GEN_2438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2440 = 7'h5e == _myNewVec_110_T_3[6:0] ? myVec_94 : _GEN_2439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2441 = 7'h5f == _myNewVec_110_T_3[6:0] ? myVec_95 : _GEN_2440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2442 = 7'h60 == _myNewVec_110_T_3[6:0] ? myVec_96 : _GEN_2441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2443 = 7'h61 == _myNewVec_110_T_3[6:0] ? myVec_97 : _GEN_2442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2444 = 7'h62 == _myNewVec_110_T_3[6:0] ? myVec_98 : _GEN_2443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2445 = 7'h63 == _myNewVec_110_T_3[6:0] ? myVec_99 : _GEN_2444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2446 = 7'h64 == _myNewVec_110_T_3[6:0] ? myVec_100 : _GEN_2445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2447 = 7'h65 == _myNewVec_110_T_3[6:0] ? myVec_101 : _GEN_2446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2448 = 7'h66 == _myNewVec_110_T_3[6:0] ? myVec_102 : _GEN_2447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2449 = 7'h67 == _myNewVec_110_T_3[6:0] ? myVec_103 : _GEN_2448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2450 = 7'h68 == _myNewVec_110_T_3[6:0] ? myVec_104 : _GEN_2449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2451 = 7'h69 == _myNewVec_110_T_3[6:0] ? myVec_105 : _GEN_2450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2452 = 7'h6a == _myNewVec_110_T_3[6:0] ? myVec_106 : _GEN_2451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2453 = 7'h6b == _myNewVec_110_T_3[6:0] ? myVec_107 : _GEN_2452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2454 = 7'h6c == _myNewVec_110_T_3[6:0] ? myVec_108 : _GEN_2453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2455 = 7'h6d == _myNewVec_110_T_3[6:0] ? myVec_109 : _GEN_2454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2456 = 7'h6e == _myNewVec_110_T_3[6:0] ? myVec_110 : _GEN_2455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2457 = 7'h6f == _myNewVec_110_T_3[6:0] ? myVec_111 : _GEN_2456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2458 = 7'h70 == _myNewVec_110_T_3[6:0] ? myVec_112 : _GEN_2457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2459 = 7'h71 == _myNewVec_110_T_3[6:0] ? myVec_113 : _GEN_2458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2460 = 7'h72 == _myNewVec_110_T_3[6:0] ? myVec_114 : _GEN_2459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2461 = 7'h73 == _myNewVec_110_T_3[6:0] ? myVec_115 : _GEN_2460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2462 = 7'h74 == _myNewVec_110_T_3[6:0] ? myVec_116 : _GEN_2461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2463 = 7'h75 == _myNewVec_110_T_3[6:0] ? myVec_117 : _GEN_2462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2464 = 7'h76 == _myNewVec_110_T_3[6:0] ? myVec_118 : _GEN_2463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2465 = 7'h77 == _myNewVec_110_T_3[6:0] ? myVec_119 : _GEN_2464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2466 = 7'h78 == _myNewVec_110_T_3[6:0] ? myVec_120 : _GEN_2465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2467 = 7'h79 == _myNewVec_110_T_3[6:0] ? myVec_121 : _GEN_2466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2468 = 7'h7a == _myNewVec_110_T_3[6:0] ? myVec_122 : _GEN_2467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2469 = 7'h7b == _myNewVec_110_T_3[6:0] ? myVec_123 : _GEN_2468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2470 = 7'h7c == _myNewVec_110_T_3[6:0] ? myVec_124 : _GEN_2469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2471 = 7'h7d == _myNewVec_110_T_3[6:0] ? myVec_125 : _GEN_2470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2472 = 7'h7e == _myNewVec_110_T_3[6:0] ? myVec_126 : _GEN_2471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_110 = 7'h7f == _myNewVec_110_T_3[6:0] ? myVec_127 : _GEN_2472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_109_T_3 = _myNewVec_127_T_1 + 16'h12; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2475 = 7'h1 == _myNewVec_109_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2476 = 7'h2 == _myNewVec_109_T_3[6:0] ? myVec_2 : _GEN_2475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2477 = 7'h3 == _myNewVec_109_T_3[6:0] ? myVec_3 : _GEN_2476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2478 = 7'h4 == _myNewVec_109_T_3[6:0] ? myVec_4 : _GEN_2477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2479 = 7'h5 == _myNewVec_109_T_3[6:0] ? myVec_5 : _GEN_2478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2480 = 7'h6 == _myNewVec_109_T_3[6:0] ? myVec_6 : _GEN_2479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2481 = 7'h7 == _myNewVec_109_T_3[6:0] ? myVec_7 : _GEN_2480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2482 = 7'h8 == _myNewVec_109_T_3[6:0] ? myVec_8 : _GEN_2481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2483 = 7'h9 == _myNewVec_109_T_3[6:0] ? myVec_9 : _GEN_2482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2484 = 7'ha == _myNewVec_109_T_3[6:0] ? myVec_10 : _GEN_2483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2485 = 7'hb == _myNewVec_109_T_3[6:0] ? myVec_11 : _GEN_2484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2486 = 7'hc == _myNewVec_109_T_3[6:0] ? myVec_12 : _GEN_2485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2487 = 7'hd == _myNewVec_109_T_3[6:0] ? myVec_13 : _GEN_2486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2488 = 7'he == _myNewVec_109_T_3[6:0] ? myVec_14 : _GEN_2487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2489 = 7'hf == _myNewVec_109_T_3[6:0] ? myVec_15 : _GEN_2488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2490 = 7'h10 == _myNewVec_109_T_3[6:0] ? myVec_16 : _GEN_2489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2491 = 7'h11 == _myNewVec_109_T_3[6:0] ? myVec_17 : _GEN_2490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2492 = 7'h12 == _myNewVec_109_T_3[6:0] ? myVec_18 : _GEN_2491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2493 = 7'h13 == _myNewVec_109_T_3[6:0] ? myVec_19 : _GEN_2492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2494 = 7'h14 == _myNewVec_109_T_3[6:0] ? myVec_20 : _GEN_2493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2495 = 7'h15 == _myNewVec_109_T_3[6:0] ? myVec_21 : _GEN_2494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2496 = 7'h16 == _myNewVec_109_T_3[6:0] ? myVec_22 : _GEN_2495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2497 = 7'h17 == _myNewVec_109_T_3[6:0] ? myVec_23 : _GEN_2496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2498 = 7'h18 == _myNewVec_109_T_3[6:0] ? myVec_24 : _GEN_2497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2499 = 7'h19 == _myNewVec_109_T_3[6:0] ? myVec_25 : _GEN_2498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2500 = 7'h1a == _myNewVec_109_T_3[6:0] ? myVec_26 : _GEN_2499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2501 = 7'h1b == _myNewVec_109_T_3[6:0] ? myVec_27 : _GEN_2500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2502 = 7'h1c == _myNewVec_109_T_3[6:0] ? myVec_28 : _GEN_2501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2503 = 7'h1d == _myNewVec_109_T_3[6:0] ? myVec_29 : _GEN_2502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2504 = 7'h1e == _myNewVec_109_T_3[6:0] ? myVec_30 : _GEN_2503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2505 = 7'h1f == _myNewVec_109_T_3[6:0] ? myVec_31 : _GEN_2504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2506 = 7'h20 == _myNewVec_109_T_3[6:0] ? myVec_32 : _GEN_2505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2507 = 7'h21 == _myNewVec_109_T_3[6:0] ? myVec_33 : _GEN_2506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2508 = 7'h22 == _myNewVec_109_T_3[6:0] ? myVec_34 : _GEN_2507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2509 = 7'h23 == _myNewVec_109_T_3[6:0] ? myVec_35 : _GEN_2508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2510 = 7'h24 == _myNewVec_109_T_3[6:0] ? myVec_36 : _GEN_2509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2511 = 7'h25 == _myNewVec_109_T_3[6:0] ? myVec_37 : _GEN_2510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2512 = 7'h26 == _myNewVec_109_T_3[6:0] ? myVec_38 : _GEN_2511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2513 = 7'h27 == _myNewVec_109_T_3[6:0] ? myVec_39 : _GEN_2512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2514 = 7'h28 == _myNewVec_109_T_3[6:0] ? myVec_40 : _GEN_2513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2515 = 7'h29 == _myNewVec_109_T_3[6:0] ? myVec_41 : _GEN_2514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2516 = 7'h2a == _myNewVec_109_T_3[6:0] ? myVec_42 : _GEN_2515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2517 = 7'h2b == _myNewVec_109_T_3[6:0] ? myVec_43 : _GEN_2516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2518 = 7'h2c == _myNewVec_109_T_3[6:0] ? myVec_44 : _GEN_2517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2519 = 7'h2d == _myNewVec_109_T_3[6:0] ? myVec_45 : _GEN_2518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2520 = 7'h2e == _myNewVec_109_T_3[6:0] ? myVec_46 : _GEN_2519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2521 = 7'h2f == _myNewVec_109_T_3[6:0] ? myVec_47 : _GEN_2520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2522 = 7'h30 == _myNewVec_109_T_3[6:0] ? myVec_48 : _GEN_2521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2523 = 7'h31 == _myNewVec_109_T_3[6:0] ? myVec_49 : _GEN_2522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2524 = 7'h32 == _myNewVec_109_T_3[6:0] ? myVec_50 : _GEN_2523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2525 = 7'h33 == _myNewVec_109_T_3[6:0] ? myVec_51 : _GEN_2524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2526 = 7'h34 == _myNewVec_109_T_3[6:0] ? myVec_52 : _GEN_2525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2527 = 7'h35 == _myNewVec_109_T_3[6:0] ? myVec_53 : _GEN_2526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2528 = 7'h36 == _myNewVec_109_T_3[6:0] ? myVec_54 : _GEN_2527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2529 = 7'h37 == _myNewVec_109_T_3[6:0] ? myVec_55 : _GEN_2528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2530 = 7'h38 == _myNewVec_109_T_3[6:0] ? myVec_56 : _GEN_2529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2531 = 7'h39 == _myNewVec_109_T_3[6:0] ? myVec_57 : _GEN_2530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2532 = 7'h3a == _myNewVec_109_T_3[6:0] ? myVec_58 : _GEN_2531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2533 = 7'h3b == _myNewVec_109_T_3[6:0] ? myVec_59 : _GEN_2532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2534 = 7'h3c == _myNewVec_109_T_3[6:0] ? myVec_60 : _GEN_2533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2535 = 7'h3d == _myNewVec_109_T_3[6:0] ? myVec_61 : _GEN_2534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2536 = 7'h3e == _myNewVec_109_T_3[6:0] ? myVec_62 : _GEN_2535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2537 = 7'h3f == _myNewVec_109_T_3[6:0] ? myVec_63 : _GEN_2536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2538 = 7'h40 == _myNewVec_109_T_3[6:0] ? myVec_64 : _GEN_2537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2539 = 7'h41 == _myNewVec_109_T_3[6:0] ? myVec_65 : _GEN_2538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2540 = 7'h42 == _myNewVec_109_T_3[6:0] ? myVec_66 : _GEN_2539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2541 = 7'h43 == _myNewVec_109_T_3[6:0] ? myVec_67 : _GEN_2540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2542 = 7'h44 == _myNewVec_109_T_3[6:0] ? myVec_68 : _GEN_2541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2543 = 7'h45 == _myNewVec_109_T_3[6:0] ? myVec_69 : _GEN_2542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2544 = 7'h46 == _myNewVec_109_T_3[6:0] ? myVec_70 : _GEN_2543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2545 = 7'h47 == _myNewVec_109_T_3[6:0] ? myVec_71 : _GEN_2544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2546 = 7'h48 == _myNewVec_109_T_3[6:0] ? myVec_72 : _GEN_2545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2547 = 7'h49 == _myNewVec_109_T_3[6:0] ? myVec_73 : _GEN_2546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2548 = 7'h4a == _myNewVec_109_T_3[6:0] ? myVec_74 : _GEN_2547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2549 = 7'h4b == _myNewVec_109_T_3[6:0] ? myVec_75 : _GEN_2548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2550 = 7'h4c == _myNewVec_109_T_3[6:0] ? myVec_76 : _GEN_2549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2551 = 7'h4d == _myNewVec_109_T_3[6:0] ? myVec_77 : _GEN_2550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2552 = 7'h4e == _myNewVec_109_T_3[6:0] ? myVec_78 : _GEN_2551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2553 = 7'h4f == _myNewVec_109_T_3[6:0] ? myVec_79 : _GEN_2552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2554 = 7'h50 == _myNewVec_109_T_3[6:0] ? myVec_80 : _GEN_2553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2555 = 7'h51 == _myNewVec_109_T_3[6:0] ? myVec_81 : _GEN_2554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2556 = 7'h52 == _myNewVec_109_T_3[6:0] ? myVec_82 : _GEN_2555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2557 = 7'h53 == _myNewVec_109_T_3[6:0] ? myVec_83 : _GEN_2556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2558 = 7'h54 == _myNewVec_109_T_3[6:0] ? myVec_84 : _GEN_2557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2559 = 7'h55 == _myNewVec_109_T_3[6:0] ? myVec_85 : _GEN_2558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2560 = 7'h56 == _myNewVec_109_T_3[6:0] ? myVec_86 : _GEN_2559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2561 = 7'h57 == _myNewVec_109_T_3[6:0] ? myVec_87 : _GEN_2560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2562 = 7'h58 == _myNewVec_109_T_3[6:0] ? myVec_88 : _GEN_2561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2563 = 7'h59 == _myNewVec_109_T_3[6:0] ? myVec_89 : _GEN_2562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2564 = 7'h5a == _myNewVec_109_T_3[6:0] ? myVec_90 : _GEN_2563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2565 = 7'h5b == _myNewVec_109_T_3[6:0] ? myVec_91 : _GEN_2564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2566 = 7'h5c == _myNewVec_109_T_3[6:0] ? myVec_92 : _GEN_2565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2567 = 7'h5d == _myNewVec_109_T_3[6:0] ? myVec_93 : _GEN_2566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2568 = 7'h5e == _myNewVec_109_T_3[6:0] ? myVec_94 : _GEN_2567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2569 = 7'h5f == _myNewVec_109_T_3[6:0] ? myVec_95 : _GEN_2568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2570 = 7'h60 == _myNewVec_109_T_3[6:0] ? myVec_96 : _GEN_2569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2571 = 7'h61 == _myNewVec_109_T_3[6:0] ? myVec_97 : _GEN_2570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2572 = 7'h62 == _myNewVec_109_T_3[6:0] ? myVec_98 : _GEN_2571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2573 = 7'h63 == _myNewVec_109_T_3[6:0] ? myVec_99 : _GEN_2572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2574 = 7'h64 == _myNewVec_109_T_3[6:0] ? myVec_100 : _GEN_2573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2575 = 7'h65 == _myNewVec_109_T_3[6:0] ? myVec_101 : _GEN_2574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2576 = 7'h66 == _myNewVec_109_T_3[6:0] ? myVec_102 : _GEN_2575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2577 = 7'h67 == _myNewVec_109_T_3[6:0] ? myVec_103 : _GEN_2576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2578 = 7'h68 == _myNewVec_109_T_3[6:0] ? myVec_104 : _GEN_2577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2579 = 7'h69 == _myNewVec_109_T_3[6:0] ? myVec_105 : _GEN_2578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2580 = 7'h6a == _myNewVec_109_T_3[6:0] ? myVec_106 : _GEN_2579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2581 = 7'h6b == _myNewVec_109_T_3[6:0] ? myVec_107 : _GEN_2580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2582 = 7'h6c == _myNewVec_109_T_3[6:0] ? myVec_108 : _GEN_2581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2583 = 7'h6d == _myNewVec_109_T_3[6:0] ? myVec_109 : _GEN_2582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2584 = 7'h6e == _myNewVec_109_T_3[6:0] ? myVec_110 : _GEN_2583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2585 = 7'h6f == _myNewVec_109_T_3[6:0] ? myVec_111 : _GEN_2584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2586 = 7'h70 == _myNewVec_109_T_3[6:0] ? myVec_112 : _GEN_2585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2587 = 7'h71 == _myNewVec_109_T_3[6:0] ? myVec_113 : _GEN_2586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2588 = 7'h72 == _myNewVec_109_T_3[6:0] ? myVec_114 : _GEN_2587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2589 = 7'h73 == _myNewVec_109_T_3[6:0] ? myVec_115 : _GEN_2588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2590 = 7'h74 == _myNewVec_109_T_3[6:0] ? myVec_116 : _GEN_2589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2591 = 7'h75 == _myNewVec_109_T_3[6:0] ? myVec_117 : _GEN_2590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2592 = 7'h76 == _myNewVec_109_T_3[6:0] ? myVec_118 : _GEN_2591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2593 = 7'h77 == _myNewVec_109_T_3[6:0] ? myVec_119 : _GEN_2592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2594 = 7'h78 == _myNewVec_109_T_3[6:0] ? myVec_120 : _GEN_2593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2595 = 7'h79 == _myNewVec_109_T_3[6:0] ? myVec_121 : _GEN_2594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2596 = 7'h7a == _myNewVec_109_T_3[6:0] ? myVec_122 : _GEN_2595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2597 = 7'h7b == _myNewVec_109_T_3[6:0] ? myVec_123 : _GEN_2596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2598 = 7'h7c == _myNewVec_109_T_3[6:0] ? myVec_124 : _GEN_2597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2599 = 7'h7d == _myNewVec_109_T_3[6:0] ? myVec_125 : _GEN_2598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2600 = 7'h7e == _myNewVec_109_T_3[6:0] ? myVec_126 : _GEN_2599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_109 = 7'h7f == _myNewVec_109_T_3[6:0] ? myVec_127 : _GEN_2600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_108_T_3 = _myNewVec_127_T_1 + 16'h13; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2603 = 7'h1 == _myNewVec_108_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2604 = 7'h2 == _myNewVec_108_T_3[6:0] ? myVec_2 : _GEN_2603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2605 = 7'h3 == _myNewVec_108_T_3[6:0] ? myVec_3 : _GEN_2604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2606 = 7'h4 == _myNewVec_108_T_3[6:0] ? myVec_4 : _GEN_2605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2607 = 7'h5 == _myNewVec_108_T_3[6:0] ? myVec_5 : _GEN_2606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2608 = 7'h6 == _myNewVec_108_T_3[6:0] ? myVec_6 : _GEN_2607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2609 = 7'h7 == _myNewVec_108_T_3[6:0] ? myVec_7 : _GEN_2608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2610 = 7'h8 == _myNewVec_108_T_3[6:0] ? myVec_8 : _GEN_2609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2611 = 7'h9 == _myNewVec_108_T_3[6:0] ? myVec_9 : _GEN_2610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2612 = 7'ha == _myNewVec_108_T_3[6:0] ? myVec_10 : _GEN_2611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2613 = 7'hb == _myNewVec_108_T_3[6:0] ? myVec_11 : _GEN_2612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2614 = 7'hc == _myNewVec_108_T_3[6:0] ? myVec_12 : _GEN_2613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2615 = 7'hd == _myNewVec_108_T_3[6:0] ? myVec_13 : _GEN_2614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2616 = 7'he == _myNewVec_108_T_3[6:0] ? myVec_14 : _GEN_2615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2617 = 7'hf == _myNewVec_108_T_3[6:0] ? myVec_15 : _GEN_2616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2618 = 7'h10 == _myNewVec_108_T_3[6:0] ? myVec_16 : _GEN_2617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2619 = 7'h11 == _myNewVec_108_T_3[6:0] ? myVec_17 : _GEN_2618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2620 = 7'h12 == _myNewVec_108_T_3[6:0] ? myVec_18 : _GEN_2619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2621 = 7'h13 == _myNewVec_108_T_3[6:0] ? myVec_19 : _GEN_2620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2622 = 7'h14 == _myNewVec_108_T_3[6:0] ? myVec_20 : _GEN_2621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2623 = 7'h15 == _myNewVec_108_T_3[6:0] ? myVec_21 : _GEN_2622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2624 = 7'h16 == _myNewVec_108_T_3[6:0] ? myVec_22 : _GEN_2623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2625 = 7'h17 == _myNewVec_108_T_3[6:0] ? myVec_23 : _GEN_2624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2626 = 7'h18 == _myNewVec_108_T_3[6:0] ? myVec_24 : _GEN_2625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2627 = 7'h19 == _myNewVec_108_T_3[6:0] ? myVec_25 : _GEN_2626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2628 = 7'h1a == _myNewVec_108_T_3[6:0] ? myVec_26 : _GEN_2627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2629 = 7'h1b == _myNewVec_108_T_3[6:0] ? myVec_27 : _GEN_2628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2630 = 7'h1c == _myNewVec_108_T_3[6:0] ? myVec_28 : _GEN_2629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2631 = 7'h1d == _myNewVec_108_T_3[6:0] ? myVec_29 : _GEN_2630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2632 = 7'h1e == _myNewVec_108_T_3[6:0] ? myVec_30 : _GEN_2631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2633 = 7'h1f == _myNewVec_108_T_3[6:0] ? myVec_31 : _GEN_2632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2634 = 7'h20 == _myNewVec_108_T_3[6:0] ? myVec_32 : _GEN_2633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2635 = 7'h21 == _myNewVec_108_T_3[6:0] ? myVec_33 : _GEN_2634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2636 = 7'h22 == _myNewVec_108_T_3[6:0] ? myVec_34 : _GEN_2635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2637 = 7'h23 == _myNewVec_108_T_3[6:0] ? myVec_35 : _GEN_2636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2638 = 7'h24 == _myNewVec_108_T_3[6:0] ? myVec_36 : _GEN_2637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2639 = 7'h25 == _myNewVec_108_T_3[6:0] ? myVec_37 : _GEN_2638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2640 = 7'h26 == _myNewVec_108_T_3[6:0] ? myVec_38 : _GEN_2639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2641 = 7'h27 == _myNewVec_108_T_3[6:0] ? myVec_39 : _GEN_2640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2642 = 7'h28 == _myNewVec_108_T_3[6:0] ? myVec_40 : _GEN_2641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2643 = 7'h29 == _myNewVec_108_T_3[6:0] ? myVec_41 : _GEN_2642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2644 = 7'h2a == _myNewVec_108_T_3[6:0] ? myVec_42 : _GEN_2643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2645 = 7'h2b == _myNewVec_108_T_3[6:0] ? myVec_43 : _GEN_2644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2646 = 7'h2c == _myNewVec_108_T_3[6:0] ? myVec_44 : _GEN_2645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2647 = 7'h2d == _myNewVec_108_T_3[6:0] ? myVec_45 : _GEN_2646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2648 = 7'h2e == _myNewVec_108_T_3[6:0] ? myVec_46 : _GEN_2647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2649 = 7'h2f == _myNewVec_108_T_3[6:0] ? myVec_47 : _GEN_2648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2650 = 7'h30 == _myNewVec_108_T_3[6:0] ? myVec_48 : _GEN_2649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2651 = 7'h31 == _myNewVec_108_T_3[6:0] ? myVec_49 : _GEN_2650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2652 = 7'h32 == _myNewVec_108_T_3[6:0] ? myVec_50 : _GEN_2651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2653 = 7'h33 == _myNewVec_108_T_3[6:0] ? myVec_51 : _GEN_2652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2654 = 7'h34 == _myNewVec_108_T_3[6:0] ? myVec_52 : _GEN_2653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2655 = 7'h35 == _myNewVec_108_T_3[6:0] ? myVec_53 : _GEN_2654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2656 = 7'h36 == _myNewVec_108_T_3[6:0] ? myVec_54 : _GEN_2655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2657 = 7'h37 == _myNewVec_108_T_3[6:0] ? myVec_55 : _GEN_2656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2658 = 7'h38 == _myNewVec_108_T_3[6:0] ? myVec_56 : _GEN_2657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2659 = 7'h39 == _myNewVec_108_T_3[6:0] ? myVec_57 : _GEN_2658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2660 = 7'h3a == _myNewVec_108_T_3[6:0] ? myVec_58 : _GEN_2659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2661 = 7'h3b == _myNewVec_108_T_3[6:0] ? myVec_59 : _GEN_2660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2662 = 7'h3c == _myNewVec_108_T_3[6:0] ? myVec_60 : _GEN_2661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2663 = 7'h3d == _myNewVec_108_T_3[6:0] ? myVec_61 : _GEN_2662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2664 = 7'h3e == _myNewVec_108_T_3[6:0] ? myVec_62 : _GEN_2663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2665 = 7'h3f == _myNewVec_108_T_3[6:0] ? myVec_63 : _GEN_2664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2666 = 7'h40 == _myNewVec_108_T_3[6:0] ? myVec_64 : _GEN_2665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2667 = 7'h41 == _myNewVec_108_T_3[6:0] ? myVec_65 : _GEN_2666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2668 = 7'h42 == _myNewVec_108_T_3[6:0] ? myVec_66 : _GEN_2667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2669 = 7'h43 == _myNewVec_108_T_3[6:0] ? myVec_67 : _GEN_2668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2670 = 7'h44 == _myNewVec_108_T_3[6:0] ? myVec_68 : _GEN_2669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2671 = 7'h45 == _myNewVec_108_T_3[6:0] ? myVec_69 : _GEN_2670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2672 = 7'h46 == _myNewVec_108_T_3[6:0] ? myVec_70 : _GEN_2671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2673 = 7'h47 == _myNewVec_108_T_3[6:0] ? myVec_71 : _GEN_2672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2674 = 7'h48 == _myNewVec_108_T_3[6:0] ? myVec_72 : _GEN_2673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2675 = 7'h49 == _myNewVec_108_T_3[6:0] ? myVec_73 : _GEN_2674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2676 = 7'h4a == _myNewVec_108_T_3[6:0] ? myVec_74 : _GEN_2675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2677 = 7'h4b == _myNewVec_108_T_3[6:0] ? myVec_75 : _GEN_2676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2678 = 7'h4c == _myNewVec_108_T_3[6:0] ? myVec_76 : _GEN_2677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2679 = 7'h4d == _myNewVec_108_T_3[6:0] ? myVec_77 : _GEN_2678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2680 = 7'h4e == _myNewVec_108_T_3[6:0] ? myVec_78 : _GEN_2679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2681 = 7'h4f == _myNewVec_108_T_3[6:0] ? myVec_79 : _GEN_2680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2682 = 7'h50 == _myNewVec_108_T_3[6:0] ? myVec_80 : _GEN_2681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2683 = 7'h51 == _myNewVec_108_T_3[6:0] ? myVec_81 : _GEN_2682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2684 = 7'h52 == _myNewVec_108_T_3[6:0] ? myVec_82 : _GEN_2683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2685 = 7'h53 == _myNewVec_108_T_3[6:0] ? myVec_83 : _GEN_2684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2686 = 7'h54 == _myNewVec_108_T_3[6:0] ? myVec_84 : _GEN_2685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2687 = 7'h55 == _myNewVec_108_T_3[6:0] ? myVec_85 : _GEN_2686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2688 = 7'h56 == _myNewVec_108_T_3[6:0] ? myVec_86 : _GEN_2687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2689 = 7'h57 == _myNewVec_108_T_3[6:0] ? myVec_87 : _GEN_2688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2690 = 7'h58 == _myNewVec_108_T_3[6:0] ? myVec_88 : _GEN_2689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2691 = 7'h59 == _myNewVec_108_T_3[6:0] ? myVec_89 : _GEN_2690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2692 = 7'h5a == _myNewVec_108_T_3[6:0] ? myVec_90 : _GEN_2691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2693 = 7'h5b == _myNewVec_108_T_3[6:0] ? myVec_91 : _GEN_2692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2694 = 7'h5c == _myNewVec_108_T_3[6:0] ? myVec_92 : _GEN_2693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2695 = 7'h5d == _myNewVec_108_T_3[6:0] ? myVec_93 : _GEN_2694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2696 = 7'h5e == _myNewVec_108_T_3[6:0] ? myVec_94 : _GEN_2695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2697 = 7'h5f == _myNewVec_108_T_3[6:0] ? myVec_95 : _GEN_2696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2698 = 7'h60 == _myNewVec_108_T_3[6:0] ? myVec_96 : _GEN_2697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2699 = 7'h61 == _myNewVec_108_T_3[6:0] ? myVec_97 : _GEN_2698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2700 = 7'h62 == _myNewVec_108_T_3[6:0] ? myVec_98 : _GEN_2699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2701 = 7'h63 == _myNewVec_108_T_3[6:0] ? myVec_99 : _GEN_2700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2702 = 7'h64 == _myNewVec_108_T_3[6:0] ? myVec_100 : _GEN_2701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2703 = 7'h65 == _myNewVec_108_T_3[6:0] ? myVec_101 : _GEN_2702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2704 = 7'h66 == _myNewVec_108_T_3[6:0] ? myVec_102 : _GEN_2703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2705 = 7'h67 == _myNewVec_108_T_3[6:0] ? myVec_103 : _GEN_2704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2706 = 7'h68 == _myNewVec_108_T_3[6:0] ? myVec_104 : _GEN_2705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2707 = 7'h69 == _myNewVec_108_T_3[6:0] ? myVec_105 : _GEN_2706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2708 = 7'h6a == _myNewVec_108_T_3[6:0] ? myVec_106 : _GEN_2707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2709 = 7'h6b == _myNewVec_108_T_3[6:0] ? myVec_107 : _GEN_2708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2710 = 7'h6c == _myNewVec_108_T_3[6:0] ? myVec_108 : _GEN_2709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2711 = 7'h6d == _myNewVec_108_T_3[6:0] ? myVec_109 : _GEN_2710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2712 = 7'h6e == _myNewVec_108_T_3[6:0] ? myVec_110 : _GEN_2711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2713 = 7'h6f == _myNewVec_108_T_3[6:0] ? myVec_111 : _GEN_2712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2714 = 7'h70 == _myNewVec_108_T_3[6:0] ? myVec_112 : _GEN_2713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2715 = 7'h71 == _myNewVec_108_T_3[6:0] ? myVec_113 : _GEN_2714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2716 = 7'h72 == _myNewVec_108_T_3[6:0] ? myVec_114 : _GEN_2715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2717 = 7'h73 == _myNewVec_108_T_3[6:0] ? myVec_115 : _GEN_2716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2718 = 7'h74 == _myNewVec_108_T_3[6:0] ? myVec_116 : _GEN_2717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2719 = 7'h75 == _myNewVec_108_T_3[6:0] ? myVec_117 : _GEN_2718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2720 = 7'h76 == _myNewVec_108_T_3[6:0] ? myVec_118 : _GEN_2719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2721 = 7'h77 == _myNewVec_108_T_3[6:0] ? myVec_119 : _GEN_2720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2722 = 7'h78 == _myNewVec_108_T_3[6:0] ? myVec_120 : _GEN_2721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2723 = 7'h79 == _myNewVec_108_T_3[6:0] ? myVec_121 : _GEN_2722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2724 = 7'h7a == _myNewVec_108_T_3[6:0] ? myVec_122 : _GEN_2723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2725 = 7'h7b == _myNewVec_108_T_3[6:0] ? myVec_123 : _GEN_2724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2726 = 7'h7c == _myNewVec_108_T_3[6:0] ? myVec_124 : _GEN_2725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2727 = 7'h7d == _myNewVec_108_T_3[6:0] ? myVec_125 : _GEN_2726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2728 = 7'h7e == _myNewVec_108_T_3[6:0] ? myVec_126 : _GEN_2727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_108 = 7'h7f == _myNewVec_108_T_3[6:0] ? myVec_127 : _GEN_2728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_107_T_3 = _myNewVec_127_T_1 + 16'h14; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2731 = 7'h1 == _myNewVec_107_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2732 = 7'h2 == _myNewVec_107_T_3[6:0] ? myVec_2 : _GEN_2731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2733 = 7'h3 == _myNewVec_107_T_3[6:0] ? myVec_3 : _GEN_2732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2734 = 7'h4 == _myNewVec_107_T_3[6:0] ? myVec_4 : _GEN_2733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2735 = 7'h5 == _myNewVec_107_T_3[6:0] ? myVec_5 : _GEN_2734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2736 = 7'h6 == _myNewVec_107_T_3[6:0] ? myVec_6 : _GEN_2735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2737 = 7'h7 == _myNewVec_107_T_3[6:0] ? myVec_7 : _GEN_2736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2738 = 7'h8 == _myNewVec_107_T_3[6:0] ? myVec_8 : _GEN_2737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2739 = 7'h9 == _myNewVec_107_T_3[6:0] ? myVec_9 : _GEN_2738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2740 = 7'ha == _myNewVec_107_T_3[6:0] ? myVec_10 : _GEN_2739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2741 = 7'hb == _myNewVec_107_T_3[6:0] ? myVec_11 : _GEN_2740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2742 = 7'hc == _myNewVec_107_T_3[6:0] ? myVec_12 : _GEN_2741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2743 = 7'hd == _myNewVec_107_T_3[6:0] ? myVec_13 : _GEN_2742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2744 = 7'he == _myNewVec_107_T_3[6:0] ? myVec_14 : _GEN_2743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2745 = 7'hf == _myNewVec_107_T_3[6:0] ? myVec_15 : _GEN_2744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2746 = 7'h10 == _myNewVec_107_T_3[6:0] ? myVec_16 : _GEN_2745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2747 = 7'h11 == _myNewVec_107_T_3[6:0] ? myVec_17 : _GEN_2746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2748 = 7'h12 == _myNewVec_107_T_3[6:0] ? myVec_18 : _GEN_2747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2749 = 7'h13 == _myNewVec_107_T_3[6:0] ? myVec_19 : _GEN_2748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2750 = 7'h14 == _myNewVec_107_T_3[6:0] ? myVec_20 : _GEN_2749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2751 = 7'h15 == _myNewVec_107_T_3[6:0] ? myVec_21 : _GEN_2750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2752 = 7'h16 == _myNewVec_107_T_3[6:0] ? myVec_22 : _GEN_2751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2753 = 7'h17 == _myNewVec_107_T_3[6:0] ? myVec_23 : _GEN_2752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2754 = 7'h18 == _myNewVec_107_T_3[6:0] ? myVec_24 : _GEN_2753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2755 = 7'h19 == _myNewVec_107_T_3[6:0] ? myVec_25 : _GEN_2754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2756 = 7'h1a == _myNewVec_107_T_3[6:0] ? myVec_26 : _GEN_2755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2757 = 7'h1b == _myNewVec_107_T_3[6:0] ? myVec_27 : _GEN_2756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2758 = 7'h1c == _myNewVec_107_T_3[6:0] ? myVec_28 : _GEN_2757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2759 = 7'h1d == _myNewVec_107_T_3[6:0] ? myVec_29 : _GEN_2758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2760 = 7'h1e == _myNewVec_107_T_3[6:0] ? myVec_30 : _GEN_2759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2761 = 7'h1f == _myNewVec_107_T_3[6:0] ? myVec_31 : _GEN_2760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2762 = 7'h20 == _myNewVec_107_T_3[6:0] ? myVec_32 : _GEN_2761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2763 = 7'h21 == _myNewVec_107_T_3[6:0] ? myVec_33 : _GEN_2762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2764 = 7'h22 == _myNewVec_107_T_3[6:0] ? myVec_34 : _GEN_2763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2765 = 7'h23 == _myNewVec_107_T_3[6:0] ? myVec_35 : _GEN_2764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2766 = 7'h24 == _myNewVec_107_T_3[6:0] ? myVec_36 : _GEN_2765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2767 = 7'h25 == _myNewVec_107_T_3[6:0] ? myVec_37 : _GEN_2766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2768 = 7'h26 == _myNewVec_107_T_3[6:0] ? myVec_38 : _GEN_2767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2769 = 7'h27 == _myNewVec_107_T_3[6:0] ? myVec_39 : _GEN_2768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2770 = 7'h28 == _myNewVec_107_T_3[6:0] ? myVec_40 : _GEN_2769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2771 = 7'h29 == _myNewVec_107_T_3[6:0] ? myVec_41 : _GEN_2770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2772 = 7'h2a == _myNewVec_107_T_3[6:0] ? myVec_42 : _GEN_2771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2773 = 7'h2b == _myNewVec_107_T_3[6:0] ? myVec_43 : _GEN_2772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2774 = 7'h2c == _myNewVec_107_T_3[6:0] ? myVec_44 : _GEN_2773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2775 = 7'h2d == _myNewVec_107_T_3[6:0] ? myVec_45 : _GEN_2774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2776 = 7'h2e == _myNewVec_107_T_3[6:0] ? myVec_46 : _GEN_2775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2777 = 7'h2f == _myNewVec_107_T_3[6:0] ? myVec_47 : _GEN_2776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2778 = 7'h30 == _myNewVec_107_T_3[6:0] ? myVec_48 : _GEN_2777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2779 = 7'h31 == _myNewVec_107_T_3[6:0] ? myVec_49 : _GEN_2778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2780 = 7'h32 == _myNewVec_107_T_3[6:0] ? myVec_50 : _GEN_2779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2781 = 7'h33 == _myNewVec_107_T_3[6:0] ? myVec_51 : _GEN_2780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2782 = 7'h34 == _myNewVec_107_T_3[6:0] ? myVec_52 : _GEN_2781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2783 = 7'h35 == _myNewVec_107_T_3[6:0] ? myVec_53 : _GEN_2782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2784 = 7'h36 == _myNewVec_107_T_3[6:0] ? myVec_54 : _GEN_2783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2785 = 7'h37 == _myNewVec_107_T_3[6:0] ? myVec_55 : _GEN_2784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2786 = 7'h38 == _myNewVec_107_T_3[6:0] ? myVec_56 : _GEN_2785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2787 = 7'h39 == _myNewVec_107_T_3[6:0] ? myVec_57 : _GEN_2786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2788 = 7'h3a == _myNewVec_107_T_3[6:0] ? myVec_58 : _GEN_2787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2789 = 7'h3b == _myNewVec_107_T_3[6:0] ? myVec_59 : _GEN_2788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2790 = 7'h3c == _myNewVec_107_T_3[6:0] ? myVec_60 : _GEN_2789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2791 = 7'h3d == _myNewVec_107_T_3[6:0] ? myVec_61 : _GEN_2790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2792 = 7'h3e == _myNewVec_107_T_3[6:0] ? myVec_62 : _GEN_2791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2793 = 7'h3f == _myNewVec_107_T_3[6:0] ? myVec_63 : _GEN_2792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2794 = 7'h40 == _myNewVec_107_T_3[6:0] ? myVec_64 : _GEN_2793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2795 = 7'h41 == _myNewVec_107_T_3[6:0] ? myVec_65 : _GEN_2794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2796 = 7'h42 == _myNewVec_107_T_3[6:0] ? myVec_66 : _GEN_2795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2797 = 7'h43 == _myNewVec_107_T_3[6:0] ? myVec_67 : _GEN_2796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2798 = 7'h44 == _myNewVec_107_T_3[6:0] ? myVec_68 : _GEN_2797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2799 = 7'h45 == _myNewVec_107_T_3[6:0] ? myVec_69 : _GEN_2798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2800 = 7'h46 == _myNewVec_107_T_3[6:0] ? myVec_70 : _GEN_2799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2801 = 7'h47 == _myNewVec_107_T_3[6:0] ? myVec_71 : _GEN_2800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2802 = 7'h48 == _myNewVec_107_T_3[6:0] ? myVec_72 : _GEN_2801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2803 = 7'h49 == _myNewVec_107_T_3[6:0] ? myVec_73 : _GEN_2802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2804 = 7'h4a == _myNewVec_107_T_3[6:0] ? myVec_74 : _GEN_2803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2805 = 7'h4b == _myNewVec_107_T_3[6:0] ? myVec_75 : _GEN_2804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2806 = 7'h4c == _myNewVec_107_T_3[6:0] ? myVec_76 : _GEN_2805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2807 = 7'h4d == _myNewVec_107_T_3[6:0] ? myVec_77 : _GEN_2806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2808 = 7'h4e == _myNewVec_107_T_3[6:0] ? myVec_78 : _GEN_2807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2809 = 7'h4f == _myNewVec_107_T_3[6:0] ? myVec_79 : _GEN_2808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2810 = 7'h50 == _myNewVec_107_T_3[6:0] ? myVec_80 : _GEN_2809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2811 = 7'h51 == _myNewVec_107_T_3[6:0] ? myVec_81 : _GEN_2810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2812 = 7'h52 == _myNewVec_107_T_3[6:0] ? myVec_82 : _GEN_2811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2813 = 7'h53 == _myNewVec_107_T_3[6:0] ? myVec_83 : _GEN_2812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2814 = 7'h54 == _myNewVec_107_T_3[6:0] ? myVec_84 : _GEN_2813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2815 = 7'h55 == _myNewVec_107_T_3[6:0] ? myVec_85 : _GEN_2814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2816 = 7'h56 == _myNewVec_107_T_3[6:0] ? myVec_86 : _GEN_2815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2817 = 7'h57 == _myNewVec_107_T_3[6:0] ? myVec_87 : _GEN_2816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2818 = 7'h58 == _myNewVec_107_T_3[6:0] ? myVec_88 : _GEN_2817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2819 = 7'h59 == _myNewVec_107_T_3[6:0] ? myVec_89 : _GEN_2818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2820 = 7'h5a == _myNewVec_107_T_3[6:0] ? myVec_90 : _GEN_2819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2821 = 7'h5b == _myNewVec_107_T_3[6:0] ? myVec_91 : _GEN_2820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2822 = 7'h5c == _myNewVec_107_T_3[6:0] ? myVec_92 : _GEN_2821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2823 = 7'h5d == _myNewVec_107_T_3[6:0] ? myVec_93 : _GEN_2822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2824 = 7'h5e == _myNewVec_107_T_3[6:0] ? myVec_94 : _GEN_2823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2825 = 7'h5f == _myNewVec_107_T_3[6:0] ? myVec_95 : _GEN_2824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2826 = 7'h60 == _myNewVec_107_T_3[6:0] ? myVec_96 : _GEN_2825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2827 = 7'h61 == _myNewVec_107_T_3[6:0] ? myVec_97 : _GEN_2826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2828 = 7'h62 == _myNewVec_107_T_3[6:0] ? myVec_98 : _GEN_2827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2829 = 7'h63 == _myNewVec_107_T_3[6:0] ? myVec_99 : _GEN_2828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2830 = 7'h64 == _myNewVec_107_T_3[6:0] ? myVec_100 : _GEN_2829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2831 = 7'h65 == _myNewVec_107_T_3[6:0] ? myVec_101 : _GEN_2830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2832 = 7'h66 == _myNewVec_107_T_3[6:0] ? myVec_102 : _GEN_2831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2833 = 7'h67 == _myNewVec_107_T_3[6:0] ? myVec_103 : _GEN_2832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2834 = 7'h68 == _myNewVec_107_T_3[6:0] ? myVec_104 : _GEN_2833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2835 = 7'h69 == _myNewVec_107_T_3[6:0] ? myVec_105 : _GEN_2834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2836 = 7'h6a == _myNewVec_107_T_3[6:0] ? myVec_106 : _GEN_2835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2837 = 7'h6b == _myNewVec_107_T_3[6:0] ? myVec_107 : _GEN_2836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2838 = 7'h6c == _myNewVec_107_T_3[6:0] ? myVec_108 : _GEN_2837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2839 = 7'h6d == _myNewVec_107_T_3[6:0] ? myVec_109 : _GEN_2838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2840 = 7'h6e == _myNewVec_107_T_3[6:0] ? myVec_110 : _GEN_2839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2841 = 7'h6f == _myNewVec_107_T_3[6:0] ? myVec_111 : _GEN_2840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2842 = 7'h70 == _myNewVec_107_T_3[6:0] ? myVec_112 : _GEN_2841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2843 = 7'h71 == _myNewVec_107_T_3[6:0] ? myVec_113 : _GEN_2842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2844 = 7'h72 == _myNewVec_107_T_3[6:0] ? myVec_114 : _GEN_2843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2845 = 7'h73 == _myNewVec_107_T_3[6:0] ? myVec_115 : _GEN_2844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2846 = 7'h74 == _myNewVec_107_T_3[6:0] ? myVec_116 : _GEN_2845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2847 = 7'h75 == _myNewVec_107_T_3[6:0] ? myVec_117 : _GEN_2846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2848 = 7'h76 == _myNewVec_107_T_3[6:0] ? myVec_118 : _GEN_2847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2849 = 7'h77 == _myNewVec_107_T_3[6:0] ? myVec_119 : _GEN_2848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2850 = 7'h78 == _myNewVec_107_T_3[6:0] ? myVec_120 : _GEN_2849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2851 = 7'h79 == _myNewVec_107_T_3[6:0] ? myVec_121 : _GEN_2850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2852 = 7'h7a == _myNewVec_107_T_3[6:0] ? myVec_122 : _GEN_2851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2853 = 7'h7b == _myNewVec_107_T_3[6:0] ? myVec_123 : _GEN_2852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2854 = 7'h7c == _myNewVec_107_T_3[6:0] ? myVec_124 : _GEN_2853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2855 = 7'h7d == _myNewVec_107_T_3[6:0] ? myVec_125 : _GEN_2854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2856 = 7'h7e == _myNewVec_107_T_3[6:0] ? myVec_126 : _GEN_2855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_107 = 7'h7f == _myNewVec_107_T_3[6:0] ? myVec_127 : _GEN_2856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_106_T_3 = _myNewVec_127_T_1 + 16'h15; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2859 = 7'h1 == _myNewVec_106_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2860 = 7'h2 == _myNewVec_106_T_3[6:0] ? myVec_2 : _GEN_2859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2861 = 7'h3 == _myNewVec_106_T_3[6:0] ? myVec_3 : _GEN_2860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2862 = 7'h4 == _myNewVec_106_T_3[6:0] ? myVec_4 : _GEN_2861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2863 = 7'h5 == _myNewVec_106_T_3[6:0] ? myVec_5 : _GEN_2862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2864 = 7'h6 == _myNewVec_106_T_3[6:0] ? myVec_6 : _GEN_2863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2865 = 7'h7 == _myNewVec_106_T_3[6:0] ? myVec_7 : _GEN_2864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2866 = 7'h8 == _myNewVec_106_T_3[6:0] ? myVec_8 : _GEN_2865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2867 = 7'h9 == _myNewVec_106_T_3[6:0] ? myVec_9 : _GEN_2866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2868 = 7'ha == _myNewVec_106_T_3[6:0] ? myVec_10 : _GEN_2867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2869 = 7'hb == _myNewVec_106_T_3[6:0] ? myVec_11 : _GEN_2868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2870 = 7'hc == _myNewVec_106_T_3[6:0] ? myVec_12 : _GEN_2869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2871 = 7'hd == _myNewVec_106_T_3[6:0] ? myVec_13 : _GEN_2870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2872 = 7'he == _myNewVec_106_T_3[6:0] ? myVec_14 : _GEN_2871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2873 = 7'hf == _myNewVec_106_T_3[6:0] ? myVec_15 : _GEN_2872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2874 = 7'h10 == _myNewVec_106_T_3[6:0] ? myVec_16 : _GEN_2873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2875 = 7'h11 == _myNewVec_106_T_3[6:0] ? myVec_17 : _GEN_2874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2876 = 7'h12 == _myNewVec_106_T_3[6:0] ? myVec_18 : _GEN_2875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2877 = 7'h13 == _myNewVec_106_T_3[6:0] ? myVec_19 : _GEN_2876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2878 = 7'h14 == _myNewVec_106_T_3[6:0] ? myVec_20 : _GEN_2877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2879 = 7'h15 == _myNewVec_106_T_3[6:0] ? myVec_21 : _GEN_2878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2880 = 7'h16 == _myNewVec_106_T_3[6:0] ? myVec_22 : _GEN_2879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2881 = 7'h17 == _myNewVec_106_T_3[6:0] ? myVec_23 : _GEN_2880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2882 = 7'h18 == _myNewVec_106_T_3[6:0] ? myVec_24 : _GEN_2881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2883 = 7'h19 == _myNewVec_106_T_3[6:0] ? myVec_25 : _GEN_2882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2884 = 7'h1a == _myNewVec_106_T_3[6:0] ? myVec_26 : _GEN_2883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2885 = 7'h1b == _myNewVec_106_T_3[6:0] ? myVec_27 : _GEN_2884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2886 = 7'h1c == _myNewVec_106_T_3[6:0] ? myVec_28 : _GEN_2885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2887 = 7'h1d == _myNewVec_106_T_3[6:0] ? myVec_29 : _GEN_2886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2888 = 7'h1e == _myNewVec_106_T_3[6:0] ? myVec_30 : _GEN_2887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2889 = 7'h1f == _myNewVec_106_T_3[6:0] ? myVec_31 : _GEN_2888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2890 = 7'h20 == _myNewVec_106_T_3[6:0] ? myVec_32 : _GEN_2889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2891 = 7'h21 == _myNewVec_106_T_3[6:0] ? myVec_33 : _GEN_2890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2892 = 7'h22 == _myNewVec_106_T_3[6:0] ? myVec_34 : _GEN_2891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2893 = 7'h23 == _myNewVec_106_T_3[6:0] ? myVec_35 : _GEN_2892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2894 = 7'h24 == _myNewVec_106_T_3[6:0] ? myVec_36 : _GEN_2893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2895 = 7'h25 == _myNewVec_106_T_3[6:0] ? myVec_37 : _GEN_2894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2896 = 7'h26 == _myNewVec_106_T_3[6:0] ? myVec_38 : _GEN_2895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2897 = 7'h27 == _myNewVec_106_T_3[6:0] ? myVec_39 : _GEN_2896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2898 = 7'h28 == _myNewVec_106_T_3[6:0] ? myVec_40 : _GEN_2897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2899 = 7'h29 == _myNewVec_106_T_3[6:0] ? myVec_41 : _GEN_2898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2900 = 7'h2a == _myNewVec_106_T_3[6:0] ? myVec_42 : _GEN_2899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2901 = 7'h2b == _myNewVec_106_T_3[6:0] ? myVec_43 : _GEN_2900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2902 = 7'h2c == _myNewVec_106_T_3[6:0] ? myVec_44 : _GEN_2901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2903 = 7'h2d == _myNewVec_106_T_3[6:0] ? myVec_45 : _GEN_2902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2904 = 7'h2e == _myNewVec_106_T_3[6:0] ? myVec_46 : _GEN_2903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2905 = 7'h2f == _myNewVec_106_T_3[6:0] ? myVec_47 : _GEN_2904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2906 = 7'h30 == _myNewVec_106_T_3[6:0] ? myVec_48 : _GEN_2905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2907 = 7'h31 == _myNewVec_106_T_3[6:0] ? myVec_49 : _GEN_2906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2908 = 7'h32 == _myNewVec_106_T_3[6:0] ? myVec_50 : _GEN_2907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2909 = 7'h33 == _myNewVec_106_T_3[6:0] ? myVec_51 : _GEN_2908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2910 = 7'h34 == _myNewVec_106_T_3[6:0] ? myVec_52 : _GEN_2909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2911 = 7'h35 == _myNewVec_106_T_3[6:0] ? myVec_53 : _GEN_2910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2912 = 7'h36 == _myNewVec_106_T_3[6:0] ? myVec_54 : _GEN_2911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2913 = 7'h37 == _myNewVec_106_T_3[6:0] ? myVec_55 : _GEN_2912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2914 = 7'h38 == _myNewVec_106_T_3[6:0] ? myVec_56 : _GEN_2913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2915 = 7'h39 == _myNewVec_106_T_3[6:0] ? myVec_57 : _GEN_2914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2916 = 7'h3a == _myNewVec_106_T_3[6:0] ? myVec_58 : _GEN_2915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2917 = 7'h3b == _myNewVec_106_T_3[6:0] ? myVec_59 : _GEN_2916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2918 = 7'h3c == _myNewVec_106_T_3[6:0] ? myVec_60 : _GEN_2917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2919 = 7'h3d == _myNewVec_106_T_3[6:0] ? myVec_61 : _GEN_2918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2920 = 7'h3e == _myNewVec_106_T_3[6:0] ? myVec_62 : _GEN_2919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2921 = 7'h3f == _myNewVec_106_T_3[6:0] ? myVec_63 : _GEN_2920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2922 = 7'h40 == _myNewVec_106_T_3[6:0] ? myVec_64 : _GEN_2921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2923 = 7'h41 == _myNewVec_106_T_3[6:0] ? myVec_65 : _GEN_2922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2924 = 7'h42 == _myNewVec_106_T_3[6:0] ? myVec_66 : _GEN_2923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2925 = 7'h43 == _myNewVec_106_T_3[6:0] ? myVec_67 : _GEN_2924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2926 = 7'h44 == _myNewVec_106_T_3[6:0] ? myVec_68 : _GEN_2925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2927 = 7'h45 == _myNewVec_106_T_3[6:0] ? myVec_69 : _GEN_2926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2928 = 7'h46 == _myNewVec_106_T_3[6:0] ? myVec_70 : _GEN_2927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2929 = 7'h47 == _myNewVec_106_T_3[6:0] ? myVec_71 : _GEN_2928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2930 = 7'h48 == _myNewVec_106_T_3[6:0] ? myVec_72 : _GEN_2929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2931 = 7'h49 == _myNewVec_106_T_3[6:0] ? myVec_73 : _GEN_2930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2932 = 7'h4a == _myNewVec_106_T_3[6:0] ? myVec_74 : _GEN_2931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2933 = 7'h4b == _myNewVec_106_T_3[6:0] ? myVec_75 : _GEN_2932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2934 = 7'h4c == _myNewVec_106_T_3[6:0] ? myVec_76 : _GEN_2933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2935 = 7'h4d == _myNewVec_106_T_3[6:0] ? myVec_77 : _GEN_2934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2936 = 7'h4e == _myNewVec_106_T_3[6:0] ? myVec_78 : _GEN_2935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2937 = 7'h4f == _myNewVec_106_T_3[6:0] ? myVec_79 : _GEN_2936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2938 = 7'h50 == _myNewVec_106_T_3[6:0] ? myVec_80 : _GEN_2937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2939 = 7'h51 == _myNewVec_106_T_3[6:0] ? myVec_81 : _GEN_2938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2940 = 7'h52 == _myNewVec_106_T_3[6:0] ? myVec_82 : _GEN_2939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2941 = 7'h53 == _myNewVec_106_T_3[6:0] ? myVec_83 : _GEN_2940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2942 = 7'h54 == _myNewVec_106_T_3[6:0] ? myVec_84 : _GEN_2941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2943 = 7'h55 == _myNewVec_106_T_3[6:0] ? myVec_85 : _GEN_2942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2944 = 7'h56 == _myNewVec_106_T_3[6:0] ? myVec_86 : _GEN_2943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2945 = 7'h57 == _myNewVec_106_T_3[6:0] ? myVec_87 : _GEN_2944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2946 = 7'h58 == _myNewVec_106_T_3[6:0] ? myVec_88 : _GEN_2945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2947 = 7'h59 == _myNewVec_106_T_3[6:0] ? myVec_89 : _GEN_2946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2948 = 7'h5a == _myNewVec_106_T_3[6:0] ? myVec_90 : _GEN_2947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2949 = 7'h5b == _myNewVec_106_T_3[6:0] ? myVec_91 : _GEN_2948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2950 = 7'h5c == _myNewVec_106_T_3[6:0] ? myVec_92 : _GEN_2949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2951 = 7'h5d == _myNewVec_106_T_3[6:0] ? myVec_93 : _GEN_2950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2952 = 7'h5e == _myNewVec_106_T_3[6:0] ? myVec_94 : _GEN_2951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2953 = 7'h5f == _myNewVec_106_T_3[6:0] ? myVec_95 : _GEN_2952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2954 = 7'h60 == _myNewVec_106_T_3[6:0] ? myVec_96 : _GEN_2953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2955 = 7'h61 == _myNewVec_106_T_3[6:0] ? myVec_97 : _GEN_2954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2956 = 7'h62 == _myNewVec_106_T_3[6:0] ? myVec_98 : _GEN_2955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2957 = 7'h63 == _myNewVec_106_T_3[6:0] ? myVec_99 : _GEN_2956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2958 = 7'h64 == _myNewVec_106_T_3[6:0] ? myVec_100 : _GEN_2957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2959 = 7'h65 == _myNewVec_106_T_3[6:0] ? myVec_101 : _GEN_2958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2960 = 7'h66 == _myNewVec_106_T_3[6:0] ? myVec_102 : _GEN_2959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2961 = 7'h67 == _myNewVec_106_T_3[6:0] ? myVec_103 : _GEN_2960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2962 = 7'h68 == _myNewVec_106_T_3[6:0] ? myVec_104 : _GEN_2961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2963 = 7'h69 == _myNewVec_106_T_3[6:0] ? myVec_105 : _GEN_2962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2964 = 7'h6a == _myNewVec_106_T_3[6:0] ? myVec_106 : _GEN_2963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2965 = 7'h6b == _myNewVec_106_T_3[6:0] ? myVec_107 : _GEN_2964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2966 = 7'h6c == _myNewVec_106_T_3[6:0] ? myVec_108 : _GEN_2965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2967 = 7'h6d == _myNewVec_106_T_3[6:0] ? myVec_109 : _GEN_2966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2968 = 7'h6e == _myNewVec_106_T_3[6:0] ? myVec_110 : _GEN_2967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2969 = 7'h6f == _myNewVec_106_T_3[6:0] ? myVec_111 : _GEN_2968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2970 = 7'h70 == _myNewVec_106_T_3[6:0] ? myVec_112 : _GEN_2969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2971 = 7'h71 == _myNewVec_106_T_3[6:0] ? myVec_113 : _GEN_2970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2972 = 7'h72 == _myNewVec_106_T_3[6:0] ? myVec_114 : _GEN_2971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2973 = 7'h73 == _myNewVec_106_T_3[6:0] ? myVec_115 : _GEN_2972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2974 = 7'h74 == _myNewVec_106_T_3[6:0] ? myVec_116 : _GEN_2973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2975 = 7'h75 == _myNewVec_106_T_3[6:0] ? myVec_117 : _GEN_2974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2976 = 7'h76 == _myNewVec_106_T_3[6:0] ? myVec_118 : _GEN_2975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2977 = 7'h77 == _myNewVec_106_T_3[6:0] ? myVec_119 : _GEN_2976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2978 = 7'h78 == _myNewVec_106_T_3[6:0] ? myVec_120 : _GEN_2977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2979 = 7'h79 == _myNewVec_106_T_3[6:0] ? myVec_121 : _GEN_2978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2980 = 7'h7a == _myNewVec_106_T_3[6:0] ? myVec_122 : _GEN_2979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2981 = 7'h7b == _myNewVec_106_T_3[6:0] ? myVec_123 : _GEN_2980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2982 = 7'h7c == _myNewVec_106_T_3[6:0] ? myVec_124 : _GEN_2981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2983 = 7'h7d == _myNewVec_106_T_3[6:0] ? myVec_125 : _GEN_2982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2984 = 7'h7e == _myNewVec_106_T_3[6:0] ? myVec_126 : _GEN_2983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_106 = 7'h7f == _myNewVec_106_T_3[6:0] ? myVec_127 : _GEN_2984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_105_T_3 = _myNewVec_127_T_1 + 16'h16; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2987 = 7'h1 == _myNewVec_105_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2988 = 7'h2 == _myNewVec_105_T_3[6:0] ? myVec_2 : _GEN_2987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2989 = 7'h3 == _myNewVec_105_T_3[6:0] ? myVec_3 : _GEN_2988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2990 = 7'h4 == _myNewVec_105_T_3[6:0] ? myVec_4 : _GEN_2989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2991 = 7'h5 == _myNewVec_105_T_3[6:0] ? myVec_5 : _GEN_2990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2992 = 7'h6 == _myNewVec_105_T_3[6:0] ? myVec_6 : _GEN_2991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2993 = 7'h7 == _myNewVec_105_T_3[6:0] ? myVec_7 : _GEN_2992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2994 = 7'h8 == _myNewVec_105_T_3[6:0] ? myVec_8 : _GEN_2993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2995 = 7'h9 == _myNewVec_105_T_3[6:0] ? myVec_9 : _GEN_2994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2996 = 7'ha == _myNewVec_105_T_3[6:0] ? myVec_10 : _GEN_2995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2997 = 7'hb == _myNewVec_105_T_3[6:0] ? myVec_11 : _GEN_2996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2998 = 7'hc == _myNewVec_105_T_3[6:0] ? myVec_12 : _GEN_2997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2999 = 7'hd == _myNewVec_105_T_3[6:0] ? myVec_13 : _GEN_2998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3000 = 7'he == _myNewVec_105_T_3[6:0] ? myVec_14 : _GEN_2999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3001 = 7'hf == _myNewVec_105_T_3[6:0] ? myVec_15 : _GEN_3000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3002 = 7'h10 == _myNewVec_105_T_3[6:0] ? myVec_16 : _GEN_3001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3003 = 7'h11 == _myNewVec_105_T_3[6:0] ? myVec_17 : _GEN_3002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3004 = 7'h12 == _myNewVec_105_T_3[6:0] ? myVec_18 : _GEN_3003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3005 = 7'h13 == _myNewVec_105_T_3[6:0] ? myVec_19 : _GEN_3004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3006 = 7'h14 == _myNewVec_105_T_3[6:0] ? myVec_20 : _GEN_3005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3007 = 7'h15 == _myNewVec_105_T_3[6:0] ? myVec_21 : _GEN_3006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3008 = 7'h16 == _myNewVec_105_T_3[6:0] ? myVec_22 : _GEN_3007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3009 = 7'h17 == _myNewVec_105_T_3[6:0] ? myVec_23 : _GEN_3008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3010 = 7'h18 == _myNewVec_105_T_3[6:0] ? myVec_24 : _GEN_3009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3011 = 7'h19 == _myNewVec_105_T_3[6:0] ? myVec_25 : _GEN_3010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3012 = 7'h1a == _myNewVec_105_T_3[6:0] ? myVec_26 : _GEN_3011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3013 = 7'h1b == _myNewVec_105_T_3[6:0] ? myVec_27 : _GEN_3012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3014 = 7'h1c == _myNewVec_105_T_3[6:0] ? myVec_28 : _GEN_3013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3015 = 7'h1d == _myNewVec_105_T_3[6:0] ? myVec_29 : _GEN_3014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3016 = 7'h1e == _myNewVec_105_T_3[6:0] ? myVec_30 : _GEN_3015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3017 = 7'h1f == _myNewVec_105_T_3[6:0] ? myVec_31 : _GEN_3016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3018 = 7'h20 == _myNewVec_105_T_3[6:0] ? myVec_32 : _GEN_3017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3019 = 7'h21 == _myNewVec_105_T_3[6:0] ? myVec_33 : _GEN_3018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3020 = 7'h22 == _myNewVec_105_T_3[6:0] ? myVec_34 : _GEN_3019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3021 = 7'h23 == _myNewVec_105_T_3[6:0] ? myVec_35 : _GEN_3020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3022 = 7'h24 == _myNewVec_105_T_3[6:0] ? myVec_36 : _GEN_3021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3023 = 7'h25 == _myNewVec_105_T_3[6:0] ? myVec_37 : _GEN_3022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3024 = 7'h26 == _myNewVec_105_T_3[6:0] ? myVec_38 : _GEN_3023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3025 = 7'h27 == _myNewVec_105_T_3[6:0] ? myVec_39 : _GEN_3024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3026 = 7'h28 == _myNewVec_105_T_3[6:0] ? myVec_40 : _GEN_3025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3027 = 7'h29 == _myNewVec_105_T_3[6:0] ? myVec_41 : _GEN_3026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3028 = 7'h2a == _myNewVec_105_T_3[6:0] ? myVec_42 : _GEN_3027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3029 = 7'h2b == _myNewVec_105_T_3[6:0] ? myVec_43 : _GEN_3028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3030 = 7'h2c == _myNewVec_105_T_3[6:0] ? myVec_44 : _GEN_3029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3031 = 7'h2d == _myNewVec_105_T_3[6:0] ? myVec_45 : _GEN_3030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3032 = 7'h2e == _myNewVec_105_T_3[6:0] ? myVec_46 : _GEN_3031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3033 = 7'h2f == _myNewVec_105_T_3[6:0] ? myVec_47 : _GEN_3032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3034 = 7'h30 == _myNewVec_105_T_3[6:0] ? myVec_48 : _GEN_3033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3035 = 7'h31 == _myNewVec_105_T_3[6:0] ? myVec_49 : _GEN_3034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3036 = 7'h32 == _myNewVec_105_T_3[6:0] ? myVec_50 : _GEN_3035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3037 = 7'h33 == _myNewVec_105_T_3[6:0] ? myVec_51 : _GEN_3036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3038 = 7'h34 == _myNewVec_105_T_3[6:0] ? myVec_52 : _GEN_3037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3039 = 7'h35 == _myNewVec_105_T_3[6:0] ? myVec_53 : _GEN_3038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3040 = 7'h36 == _myNewVec_105_T_3[6:0] ? myVec_54 : _GEN_3039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3041 = 7'h37 == _myNewVec_105_T_3[6:0] ? myVec_55 : _GEN_3040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3042 = 7'h38 == _myNewVec_105_T_3[6:0] ? myVec_56 : _GEN_3041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3043 = 7'h39 == _myNewVec_105_T_3[6:0] ? myVec_57 : _GEN_3042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3044 = 7'h3a == _myNewVec_105_T_3[6:0] ? myVec_58 : _GEN_3043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3045 = 7'h3b == _myNewVec_105_T_3[6:0] ? myVec_59 : _GEN_3044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3046 = 7'h3c == _myNewVec_105_T_3[6:0] ? myVec_60 : _GEN_3045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3047 = 7'h3d == _myNewVec_105_T_3[6:0] ? myVec_61 : _GEN_3046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3048 = 7'h3e == _myNewVec_105_T_3[6:0] ? myVec_62 : _GEN_3047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3049 = 7'h3f == _myNewVec_105_T_3[6:0] ? myVec_63 : _GEN_3048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3050 = 7'h40 == _myNewVec_105_T_3[6:0] ? myVec_64 : _GEN_3049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3051 = 7'h41 == _myNewVec_105_T_3[6:0] ? myVec_65 : _GEN_3050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3052 = 7'h42 == _myNewVec_105_T_3[6:0] ? myVec_66 : _GEN_3051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3053 = 7'h43 == _myNewVec_105_T_3[6:0] ? myVec_67 : _GEN_3052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3054 = 7'h44 == _myNewVec_105_T_3[6:0] ? myVec_68 : _GEN_3053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3055 = 7'h45 == _myNewVec_105_T_3[6:0] ? myVec_69 : _GEN_3054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3056 = 7'h46 == _myNewVec_105_T_3[6:0] ? myVec_70 : _GEN_3055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3057 = 7'h47 == _myNewVec_105_T_3[6:0] ? myVec_71 : _GEN_3056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3058 = 7'h48 == _myNewVec_105_T_3[6:0] ? myVec_72 : _GEN_3057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3059 = 7'h49 == _myNewVec_105_T_3[6:0] ? myVec_73 : _GEN_3058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3060 = 7'h4a == _myNewVec_105_T_3[6:0] ? myVec_74 : _GEN_3059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3061 = 7'h4b == _myNewVec_105_T_3[6:0] ? myVec_75 : _GEN_3060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3062 = 7'h4c == _myNewVec_105_T_3[6:0] ? myVec_76 : _GEN_3061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3063 = 7'h4d == _myNewVec_105_T_3[6:0] ? myVec_77 : _GEN_3062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3064 = 7'h4e == _myNewVec_105_T_3[6:0] ? myVec_78 : _GEN_3063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3065 = 7'h4f == _myNewVec_105_T_3[6:0] ? myVec_79 : _GEN_3064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3066 = 7'h50 == _myNewVec_105_T_3[6:0] ? myVec_80 : _GEN_3065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3067 = 7'h51 == _myNewVec_105_T_3[6:0] ? myVec_81 : _GEN_3066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3068 = 7'h52 == _myNewVec_105_T_3[6:0] ? myVec_82 : _GEN_3067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3069 = 7'h53 == _myNewVec_105_T_3[6:0] ? myVec_83 : _GEN_3068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3070 = 7'h54 == _myNewVec_105_T_3[6:0] ? myVec_84 : _GEN_3069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3071 = 7'h55 == _myNewVec_105_T_3[6:0] ? myVec_85 : _GEN_3070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3072 = 7'h56 == _myNewVec_105_T_3[6:0] ? myVec_86 : _GEN_3071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3073 = 7'h57 == _myNewVec_105_T_3[6:0] ? myVec_87 : _GEN_3072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3074 = 7'h58 == _myNewVec_105_T_3[6:0] ? myVec_88 : _GEN_3073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3075 = 7'h59 == _myNewVec_105_T_3[6:0] ? myVec_89 : _GEN_3074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3076 = 7'h5a == _myNewVec_105_T_3[6:0] ? myVec_90 : _GEN_3075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3077 = 7'h5b == _myNewVec_105_T_3[6:0] ? myVec_91 : _GEN_3076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3078 = 7'h5c == _myNewVec_105_T_3[6:0] ? myVec_92 : _GEN_3077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3079 = 7'h5d == _myNewVec_105_T_3[6:0] ? myVec_93 : _GEN_3078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3080 = 7'h5e == _myNewVec_105_T_3[6:0] ? myVec_94 : _GEN_3079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3081 = 7'h5f == _myNewVec_105_T_3[6:0] ? myVec_95 : _GEN_3080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3082 = 7'h60 == _myNewVec_105_T_3[6:0] ? myVec_96 : _GEN_3081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3083 = 7'h61 == _myNewVec_105_T_3[6:0] ? myVec_97 : _GEN_3082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3084 = 7'h62 == _myNewVec_105_T_3[6:0] ? myVec_98 : _GEN_3083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3085 = 7'h63 == _myNewVec_105_T_3[6:0] ? myVec_99 : _GEN_3084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3086 = 7'h64 == _myNewVec_105_T_3[6:0] ? myVec_100 : _GEN_3085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3087 = 7'h65 == _myNewVec_105_T_3[6:0] ? myVec_101 : _GEN_3086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3088 = 7'h66 == _myNewVec_105_T_3[6:0] ? myVec_102 : _GEN_3087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3089 = 7'h67 == _myNewVec_105_T_3[6:0] ? myVec_103 : _GEN_3088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3090 = 7'h68 == _myNewVec_105_T_3[6:0] ? myVec_104 : _GEN_3089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3091 = 7'h69 == _myNewVec_105_T_3[6:0] ? myVec_105 : _GEN_3090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3092 = 7'h6a == _myNewVec_105_T_3[6:0] ? myVec_106 : _GEN_3091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3093 = 7'h6b == _myNewVec_105_T_3[6:0] ? myVec_107 : _GEN_3092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3094 = 7'h6c == _myNewVec_105_T_3[6:0] ? myVec_108 : _GEN_3093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3095 = 7'h6d == _myNewVec_105_T_3[6:0] ? myVec_109 : _GEN_3094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3096 = 7'h6e == _myNewVec_105_T_3[6:0] ? myVec_110 : _GEN_3095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3097 = 7'h6f == _myNewVec_105_T_3[6:0] ? myVec_111 : _GEN_3096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3098 = 7'h70 == _myNewVec_105_T_3[6:0] ? myVec_112 : _GEN_3097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3099 = 7'h71 == _myNewVec_105_T_3[6:0] ? myVec_113 : _GEN_3098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3100 = 7'h72 == _myNewVec_105_T_3[6:0] ? myVec_114 : _GEN_3099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3101 = 7'h73 == _myNewVec_105_T_3[6:0] ? myVec_115 : _GEN_3100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3102 = 7'h74 == _myNewVec_105_T_3[6:0] ? myVec_116 : _GEN_3101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3103 = 7'h75 == _myNewVec_105_T_3[6:0] ? myVec_117 : _GEN_3102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3104 = 7'h76 == _myNewVec_105_T_3[6:0] ? myVec_118 : _GEN_3103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3105 = 7'h77 == _myNewVec_105_T_3[6:0] ? myVec_119 : _GEN_3104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3106 = 7'h78 == _myNewVec_105_T_3[6:0] ? myVec_120 : _GEN_3105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3107 = 7'h79 == _myNewVec_105_T_3[6:0] ? myVec_121 : _GEN_3106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3108 = 7'h7a == _myNewVec_105_T_3[6:0] ? myVec_122 : _GEN_3107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3109 = 7'h7b == _myNewVec_105_T_3[6:0] ? myVec_123 : _GEN_3108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3110 = 7'h7c == _myNewVec_105_T_3[6:0] ? myVec_124 : _GEN_3109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3111 = 7'h7d == _myNewVec_105_T_3[6:0] ? myVec_125 : _GEN_3110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3112 = 7'h7e == _myNewVec_105_T_3[6:0] ? myVec_126 : _GEN_3111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_105 = 7'h7f == _myNewVec_105_T_3[6:0] ? myVec_127 : _GEN_3112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_104_T_3 = _myNewVec_127_T_1 + 16'h17; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3115 = 7'h1 == _myNewVec_104_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3116 = 7'h2 == _myNewVec_104_T_3[6:0] ? myVec_2 : _GEN_3115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3117 = 7'h3 == _myNewVec_104_T_3[6:0] ? myVec_3 : _GEN_3116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3118 = 7'h4 == _myNewVec_104_T_3[6:0] ? myVec_4 : _GEN_3117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3119 = 7'h5 == _myNewVec_104_T_3[6:0] ? myVec_5 : _GEN_3118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3120 = 7'h6 == _myNewVec_104_T_3[6:0] ? myVec_6 : _GEN_3119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3121 = 7'h7 == _myNewVec_104_T_3[6:0] ? myVec_7 : _GEN_3120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3122 = 7'h8 == _myNewVec_104_T_3[6:0] ? myVec_8 : _GEN_3121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3123 = 7'h9 == _myNewVec_104_T_3[6:0] ? myVec_9 : _GEN_3122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3124 = 7'ha == _myNewVec_104_T_3[6:0] ? myVec_10 : _GEN_3123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3125 = 7'hb == _myNewVec_104_T_3[6:0] ? myVec_11 : _GEN_3124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3126 = 7'hc == _myNewVec_104_T_3[6:0] ? myVec_12 : _GEN_3125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3127 = 7'hd == _myNewVec_104_T_3[6:0] ? myVec_13 : _GEN_3126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3128 = 7'he == _myNewVec_104_T_3[6:0] ? myVec_14 : _GEN_3127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3129 = 7'hf == _myNewVec_104_T_3[6:0] ? myVec_15 : _GEN_3128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3130 = 7'h10 == _myNewVec_104_T_3[6:0] ? myVec_16 : _GEN_3129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3131 = 7'h11 == _myNewVec_104_T_3[6:0] ? myVec_17 : _GEN_3130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3132 = 7'h12 == _myNewVec_104_T_3[6:0] ? myVec_18 : _GEN_3131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3133 = 7'h13 == _myNewVec_104_T_3[6:0] ? myVec_19 : _GEN_3132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3134 = 7'h14 == _myNewVec_104_T_3[6:0] ? myVec_20 : _GEN_3133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3135 = 7'h15 == _myNewVec_104_T_3[6:0] ? myVec_21 : _GEN_3134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3136 = 7'h16 == _myNewVec_104_T_3[6:0] ? myVec_22 : _GEN_3135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3137 = 7'h17 == _myNewVec_104_T_3[6:0] ? myVec_23 : _GEN_3136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3138 = 7'h18 == _myNewVec_104_T_3[6:0] ? myVec_24 : _GEN_3137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3139 = 7'h19 == _myNewVec_104_T_3[6:0] ? myVec_25 : _GEN_3138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3140 = 7'h1a == _myNewVec_104_T_3[6:0] ? myVec_26 : _GEN_3139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3141 = 7'h1b == _myNewVec_104_T_3[6:0] ? myVec_27 : _GEN_3140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3142 = 7'h1c == _myNewVec_104_T_3[6:0] ? myVec_28 : _GEN_3141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3143 = 7'h1d == _myNewVec_104_T_3[6:0] ? myVec_29 : _GEN_3142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3144 = 7'h1e == _myNewVec_104_T_3[6:0] ? myVec_30 : _GEN_3143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3145 = 7'h1f == _myNewVec_104_T_3[6:0] ? myVec_31 : _GEN_3144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3146 = 7'h20 == _myNewVec_104_T_3[6:0] ? myVec_32 : _GEN_3145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3147 = 7'h21 == _myNewVec_104_T_3[6:0] ? myVec_33 : _GEN_3146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3148 = 7'h22 == _myNewVec_104_T_3[6:0] ? myVec_34 : _GEN_3147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3149 = 7'h23 == _myNewVec_104_T_3[6:0] ? myVec_35 : _GEN_3148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3150 = 7'h24 == _myNewVec_104_T_3[6:0] ? myVec_36 : _GEN_3149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3151 = 7'h25 == _myNewVec_104_T_3[6:0] ? myVec_37 : _GEN_3150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3152 = 7'h26 == _myNewVec_104_T_3[6:0] ? myVec_38 : _GEN_3151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3153 = 7'h27 == _myNewVec_104_T_3[6:0] ? myVec_39 : _GEN_3152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3154 = 7'h28 == _myNewVec_104_T_3[6:0] ? myVec_40 : _GEN_3153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3155 = 7'h29 == _myNewVec_104_T_3[6:0] ? myVec_41 : _GEN_3154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3156 = 7'h2a == _myNewVec_104_T_3[6:0] ? myVec_42 : _GEN_3155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3157 = 7'h2b == _myNewVec_104_T_3[6:0] ? myVec_43 : _GEN_3156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3158 = 7'h2c == _myNewVec_104_T_3[6:0] ? myVec_44 : _GEN_3157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3159 = 7'h2d == _myNewVec_104_T_3[6:0] ? myVec_45 : _GEN_3158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3160 = 7'h2e == _myNewVec_104_T_3[6:0] ? myVec_46 : _GEN_3159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3161 = 7'h2f == _myNewVec_104_T_3[6:0] ? myVec_47 : _GEN_3160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3162 = 7'h30 == _myNewVec_104_T_3[6:0] ? myVec_48 : _GEN_3161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3163 = 7'h31 == _myNewVec_104_T_3[6:0] ? myVec_49 : _GEN_3162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3164 = 7'h32 == _myNewVec_104_T_3[6:0] ? myVec_50 : _GEN_3163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3165 = 7'h33 == _myNewVec_104_T_3[6:0] ? myVec_51 : _GEN_3164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3166 = 7'h34 == _myNewVec_104_T_3[6:0] ? myVec_52 : _GEN_3165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3167 = 7'h35 == _myNewVec_104_T_3[6:0] ? myVec_53 : _GEN_3166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3168 = 7'h36 == _myNewVec_104_T_3[6:0] ? myVec_54 : _GEN_3167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3169 = 7'h37 == _myNewVec_104_T_3[6:0] ? myVec_55 : _GEN_3168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3170 = 7'h38 == _myNewVec_104_T_3[6:0] ? myVec_56 : _GEN_3169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3171 = 7'h39 == _myNewVec_104_T_3[6:0] ? myVec_57 : _GEN_3170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3172 = 7'h3a == _myNewVec_104_T_3[6:0] ? myVec_58 : _GEN_3171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3173 = 7'h3b == _myNewVec_104_T_3[6:0] ? myVec_59 : _GEN_3172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3174 = 7'h3c == _myNewVec_104_T_3[6:0] ? myVec_60 : _GEN_3173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3175 = 7'h3d == _myNewVec_104_T_3[6:0] ? myVec_61 : _GEN_3174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3176 = 7'h3e == _myNewVec_104_T_3[6:0] ? myVec_62 : _GEN_3175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3177 = 7'h3f == _myNewVec_104_T_3[6:0] ? myVec_63 : _GEN_3176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3178 = 7'h40 == _myNewVec_104_T_3[6:0] ? myVec_64 : _GEN_3177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3179 = 7'h41 == _myNewVec_104_T_3[6:0] ? myVec_65 : _GEN_3178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3180 = 7'h42 == _myNewVec_104_T_3[6:0] ? myVec_66 : _GEN_3179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3181 = 7'h43 == _myNewVec_104_T_3[6:0] ? myVec_67 : _GEN_3180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3182 = 7'h44 == _myNewVec_104_T_3[6:0] ? myVec_68 : _GEN_3181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3183 = 7'h45 == _myNewVec_104_T_3[6:0] ? myVec_69 : _GEN_3182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3184 = 7'h46 == _myNewVec_104_T_3[6:0] ? myVec_70 : _GEN_3183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3185 = 7'h47 == _myNewVec_104_T_3[6:0] ? myVec_71 : _GEN_3184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3186 = 7'h48 == _myNewVec_104_T_3[6:0] ? myVec_72 : _GEN_3185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3187 = 7'h49 == _myNewVec_104_T_3[6:0] ? myVec_73 : _GEN_3186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3188 = 7'h4a == _myNewVec_104_T_3[6:0] ? myVec_74 : _GEN_3187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3189 = 7'h4b == _myNewVec_104_T_3[6:0] ? myVec_75 : _GEN_3188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3190 = 7'h4c == _myNewVec_104_T_3[6:0] ? myVec_76 : _GEN_3189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3191 = 7'h4d == _myNewVec_104_T_3[6:0] ? myVec_77 : _GEN_3190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3192 = 7'h4e == _myNewVec_104_T_3[6:0] ? myVec_78 : _GEN_3191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3193 = 7'h4f == _myNewVec_104_T_3[6:0] ? myVec_79 : _GEN_3192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3194 = 7'h50 == _myNewVec_104_T_3[6:0] ? myVec_80 : _GEN_3193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3195 = 7'h51 == _myNewVec_104_T_3[6:0] ? myVec_81 : _GEN_3194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3196 = 7'h52 == _myNewVec_104_T_3[6:0] ? myVec_82 : _GEN_3195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3197 = 7'h53 == _myNewVec_104_T_3[6:0] ? myVec_83 : _GEN_3196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3198 = 7'h54 == _myNewVec_104_T_3[6:0] ? myVec_84 : _GEN_3197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3199 = 7'h55 == _myNewVec_104_T_3[6:0] ? myVec_85 : _GEN_3198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3200 = 7'h56 == _myNewVec_104_T_3[6:0] ? myVec_86 : _GEN_3199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3201 = 7'h57 == _myNewVec_104_T_3[6:0] ? myVec_87 : _GEN_3200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3202 = 7'h58 == _myNewVec_104_T_3[6:0] ? myVec_88 : _GEN_3201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3203 = 7'h59 == _myNewVec_104_T_3[6:0] ? myVec_89 : _GEN_3202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3204 = 7'h5a == _myNewVec_104_T_3[6:0] ? myVec_90 : _GEN_3203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3205 = 7'h5b == _myNewVec_104_T_3[6:0] ? myVec_91 : _GEN_3204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3206 = 7'h5c == _myNewVec_104_T_3[6:0] ? myVec_92 : _GEN_3205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3207 = 7'h5d == _myNewVec_104_T_3[6:0] ? myVec_93 : _GEN_3206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3208 = 7'h5e == _myNewVec_104_T_3[6:0] ? myVec_94 : _GEN_3207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3209 = 7'h5f == _myNewVec_104_T_3[6:0] ? myVec_95 : _GEN_3208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3210 = 7'h60 == _myNewVec_104_T_3[6:0] ? myVec_96 : _GEN_3209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3211 = 7'h61 == _myNewVec_104_T_3[6:0] ? myVec_97 : _GEN_3210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3212 = 7'h62 == _myNewVec_104_T_3[6:0] ? myVec_98 : _GEN_3211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3213 = 7'h63 == _myNewVec_104_T_3[6:0] ? myVec_99 : _GEN_3212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3214 = 7'h64 == _myNewVec_104_T_3[6:0] ? myVec_100 : _GEN_3213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3215 = 7'h65 == _myNewVec_104_T_3[6:0] ? myVec_101 : _GEN_3214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3216 = 7'h66 == _myNewVec_104_T_3[6:0] ? myVec_102 : _GEN_3215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3217 = 7'h67 == _myNewVec_104_T_3[6:0] ? myVec_103 : _GEN_3216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3218 = 7'h68 == _myNewVec_104_T_3[6:0] ? myVec_104 : _GEN_3217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3219 = 7'h69 == _myNewVec_104_T_3[6:0] ? myVec_105 : _GEN_3218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3220 = 7'h6a == _myNewVec_104_T_3[6:0] ? myVec_106 : _GEN_3219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3221 = 7'h6b == _myNewVec_104_T_3[6:0] ? myVec_107 : _GEN_3220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3222 = 7'h6c == _myNewVec_104_T_3[6:0] ? myVec_108 : _GEN_3221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3223 = 7'h6d == _myNewVec_104_T_3[6:0] ? myVec_109 : _GEN_3222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3224 = 7'h6e == _myNewVec_104_T_3[6:0] ? myVec_110 : _GEN_3223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3225 = 7'h6f == _myNewVec_104_T_3[6:0] ? myVec_111 : _GEN_3224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3226 = 7'h70 == _myNewVec_104_T_3[6:0] ? myVec_112 : _GEN_3225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3227 = 7'h71 == _myNewVec_104_T_3[6:0] ? myVec_113 : _GEN_3226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3228 = 7'h72 == _myNewVec_104_T_3[6:0] ? myVec_114 : _GEN_3227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3229 = 7'h73 == _myNewVec_104_T_3[6:0] ? myVec_115 : _GEN_3228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3230 = 7'h74 == _myNewVec_104_T_3[6:0] ? myVec_116 : _GEN_3229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3231 = 7'h75 == _myNewVec_104_T_3[6:0] ? myVec_117 : _GEN_3230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3232 = 7'h76 == _myNewVec_104_T_3[6:0] ? myVec_118 : _GEN_3231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3233 = 7'h77 == _myNewVec_104_T_3[6:0] ? myVec_119 : _GEN_3232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3234 = 7'h78 == _myNewVec_104_T_3[6:0] ? myVec_120 : _GEN_3233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3235 = 7'h79 == _myNewVec_104_T_3[6:0] ? myVec_121 : _GEN_3234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3236 = 7'h7a == _myNewVec_104_T_3[6:0] ? myVec_122 : _GEN_3235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3237 = 7'h7b == _myNewVec_104_T_3[6:0] ? myVec_123 : _GEN_3236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3238 = 7'h7c == _myNewVec_104_T_3[6:0] ? myVec_124 : _GEN_3237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3239 = 7'h7d == _myNewVec_104_T_3[6:0] ? myVec_125 : _GEN_3238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3240 = 7'h7e == _myNewVec_104_T_3[6:0] ? myVec_126 : _GEN_3239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_104 = 7'h7f == _myNewVec_104_T_3[6:0] ? myVec_127 : _GEN_3240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_103_T_3 = _myNewVec_127_T_1 + 16'h18; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3243 = 7'h1 == _myNewVec_103_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3244 = 7'h2 == _myNewVec_103_T_3[6:0] ? myVec_2 : _GEN_3243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3245 = 7'h3 == _myNewVec_103_T_3[6:0] ? myVec_3 : _GEN_3244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3246 = 7'h4 == _myNewVec_103_T_3[6:0] ? myVec_4 : _GEN_3245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3247 = 7'h5 == _myNewVec_103_T_3[6:0] ? myVec_5 : _GEN_3246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3248 = 7'h6 == _myNewVec_103_T_3[6:0] ? myVec_6 : _GEN_3247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3249 = 7'h7 == _myNewVec_103_T_3[6:0] ? myVec_7 : _GEN_3248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3250 = 7'h8 == _myNewVec_103_T_3[6:0] ? myVec_8 : _GEN_3249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3251 = 7'h9 == _myNewVec_103_T_3[6:0] ? myVec_9 : _GEN_3250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3252 = 7'ha == _myNewVec_103_T_3[6:0] ? myVec_10 : _GEN_3251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3253 = 7'hb == _myNewVec_103_T_3[6:0] ? myVec_11 : _GEN_3252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3254 = 7'hc == _myNewVec_103_T_3[6:0] ? myVec_12 : _GEN_3253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3255 = 7'hd == _myNewVec_103_T_3[6:0] ? myVec_13 : _GEN_3254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3256 = 7'he == _myNewVec_103_T_3[6:0] ? myVec_14 : _GEN_3255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3257 = 7'hf == _myNewVec_103_T_3[6:0] ? myVec_15 : _GEN_3256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3258 = 7'h10 == _myNewVec_103_T_3[6:0] ? myVec_16 : _GEN_3257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3259 = 7'h11 == _myNewVec_103_T_3[6:0] ? myVec_17 : _GEN_3258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3260 = 7'h12 == _myNewVec_103_T_3[6:0] ? myVec_18 : _GEN_3259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3261 = 7'h13 == _myNewVec_103_T_3[6:0] ? myVec_19 : _GEN_3260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3262 = 7'h14 == _myNewVec_103_T_3[6:0] ? myVec_20 : _GEN_3261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3263 = 7'h15 == _myNewVec_103_T_3[6:0] ? myVec_21 : _GEN_3262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3264 = 7'h16 == _myNewVec_103_T_3[6:0] ? myVec_22 : _GEN_3263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3265 = 7'h17 == _myNewVec_103_T_3[6:0] ? myVec_23 : _GEN_3264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3266 = 7'h18 == _myNewVec_103_T_3[6:0] ? myVec_24 : _GEN_3265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3267 = 7'h19 == _myNewVec_103_T_3[6:0] ? myVec_25 : _GEN_3266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3268 = 7'h1a == _myNewVec_103_T_3[6:0] ? myVec_26 : _GEN_3267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3269 = 7'h1b == _myNewVec_103_T_3[6:0] ? myVec_27 : _GEN_3268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3270 = 7'h1c == _myNewVec_103_T_3[6:0] ? myVec_28 : _GEN_3269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3271 = 7'h1d == _myNewVec_103_T_3[6:0] ? myVec_29 : _GEN_3270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3272 = 7'h1e == _myNewVec_103_T_3[6:0] ? myVec_30 : _GEN_3271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3273 = 7'h1f == _myNewVec_103_T_3[6:0] ? myVec_31 : _GEN_3272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3274 = 7'h20 == _myNewVec_103_T_3[6:0] ? myVec_32 : _GEN_3273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3275 = 7'h21 == _myNewVec_103_T_3[6:0] ? myVec_33 : _GEN_3274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3276 = 7'h22 == _myNewVec_103_T_3[6:0] ? myVec_34 : _GEN_3275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3277 = 7'h23 == _myNewVec_103_T_3[6:0] ? myVec_35 : _GEN_3276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3278 = 7'h24 == _myNewVec_103_T_3[6:0] ? myVec_36 : _GEN_3277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3279 = 7'h25 == _myNewVec_103_T_3[6:0] ? myVec_37 : _GEN_3278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3280 = 7'h26 == _myNewVec_103_T_3[6:0] ? myVec_38 : _GEN_3279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3281 = 7'h27 == _myNewVec_103_T_3[6:0] ? myVec_39 : _GEN_3280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3282 = 7'h28 == _myNewVec_103_T_3[6:0] ? myVec_40 : _GEN_3281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3283 = 7'h29 == _myNewVec_103_T_3[6:0] ? myVec_41 : _GEN_3282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3284 = 7'h2a == _myNewVec_103_T_3[6:0] ? myVec_42 : _GEN_3283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3285 = 7'h2b == _myNewVec_103_T_3[6:0] ? myVec_43 : _GEN_3284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3286 = 7'h2c == _myNewVec_103_T_3[6:0] ? myVec_44 : _GEN_3285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3287 = 7'h2d == _myNewVec_103_T_3[6:0] ? myVec_45 : _GEN_3286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3288 = 7'h2e == _myNewVec_103_T_3[6:0] ? myVec_46 : _GEN_3287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3289 = 7'h2f == _myNewVec_103_T_3[6:0] ? myVec_47 : _GEN_3288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3290 = 7'h30 == _myNewVec_103_T_3[6:0] ? myVec_48 : _GEN_3289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3291 = 7'h31 == _myNewVec_103_T_3[6:0] ? myVec_49 : _GEN_3290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3292 = 7'h32 == _myNewVec_103_T_3[6:0] ? myVec_50 : _GEN_3291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3293 = 7'h33 == _myNewVec_103_T_3[6:0] ? myVec_51 : _GEN_3292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3294 = 7'h34 == _myNewVec_103_T_3[6:0] ? myVec_52 : _GEN_3293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3295 = 7'h35 == _myNewVec_103_T_3[6:0] ? myVec_53 : _GEN_3294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3296 = 7'h36 == _myNewVec_103_T_3[6:0] ? myVec_54 : _GEN_3295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3297 = 7'h37 == _myNewVec_103_T_3[6:0] ? myVec_55 : _GEN_3296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3298 = 7'h38 == _myNewVec_103_T_3[6:0] ? myVec_56 : _GEN_3297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3299 = 7'h39 == _myNewVec_103_T_3[6:0] ? myVec_57 : _GEN_3298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3300 = 7'h3a == _myNewVec_103_T_3[6:0] ? myVec_58 : _GEN_3299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3301 = 7'h3b == _myNewVec_103_T_3[6:0] ? myVec_59 : _GEN_3300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3302 = 7'h3c == _myNewVec_103_T_3[6:0] ? myVec_60 : _GEN_3301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3303 = 7'h3d == _myNewVec_103_T_3[6:0] ? myVec_61 : _GEN_3302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3304 = 7'h3e == _myNewVec_103_T_3[6:0] ? myVec_62 : _GEN_3303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3305 = 7'h3f == _myNewVec_103_T_3[6:0] ? myVec_63 : _GEN_3304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3306 = 7'h40 == _myNewVec_103_T_3[6:0] ? myVec_64 : _GEN_3305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3307 = 7'h41 == _myNewVec_103_T_3[6:0] ? myVec_65 : _GEN_3306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3308 = 7'h42 == _myNewVec_103_T_3[6:0] ? myVec_66 : _GEN_3307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3309 = 7'h43 == _myNewVec_103_T_3[6:0] ? myVec_67 : _GEN_3308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3310 = 7'h44 == _myNewVec_103_T_3[6:0] ? myVec_68 : _GEN_3309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3311 = 7'h45 == _myNewVec_103_T_3[6:0] ? myVec_69 : _GEN_3310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3312 = 7'h46 == _myNewVec_103_T_3[6:0] ? myVec_70 : _GEN_3311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3313 = 7'h47 == _myNewVec_103_T_3[6:0] ? myVec_71 : _GEN_3312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3314 = 7'h48 == _myNewVec_103_T_3[6:0] ? myVec_72 : _GEN_3313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3315 = 7'h49 == _myNewVec_103_T_3[6:0] ? myVec_73 : _GEN_3314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3316 = 7'h4a == _myNewVec_103_T_3[6:0] ? myVec_74 : _GEN_3315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3317 = 7'h4b == _myNewVec_103_T_3[6:0] ? myVec_75 : _GEN_3316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3318 = 7'h4c == _myNewVec_103_T_3[6:0] ? myVec_76 : _GEN_3317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3319 = 7'h4d == _myNewVec_103_T_3[6:0] ? myVec_77 : _GEN_3318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3320 = 7'h4e == _myNewVec_103_T_3[6:0] ? myVec_78 : _GEN_3319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3321 = 7'h4f == _myNewVec_103_T_3[6:0] ? myVec_79 : _GEN_3320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3322 = 7'h50 == _myNewVec_103_T_3[6:0] ? myVec_80 : _GEN_3321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3323 = 7'h51 == _myNewVec_103_T_3[6:0] ? myVec_81 : _GEN_3322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3324 = 7'h52 == _myNewVec_103_T_3[6:0] ? myVec_82 : _GEN_3323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3325 = 7'h53 == _myNewVec_103_T_3[6:0] ? myVec_83 : _GEN_3324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3326 = 7'h54 == _myNewVec_103_T_3[6:0] ? myVec_84 : _GEN_3325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3327 = 7'h55 == _myNewVec_103_T_3[6:0] ? myVec_85 : _GEN_3326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3328 = 7'h56 == _myNewVec_103_T_3[6:0] ? myVec_86 : _GEN_3327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3329 = 7'h57 == _myNewVec_103_T_3[6:0] ? myVec_87 : _GEN_3328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3330 = 7'h58 == _myNewVec_103_T_3[6:0] ? myVec_88 : _GEN_3329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3331 = 7'h59 == _myNewVec_103_T_3[6:0] ? myVec_89 : _GEN_3330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3332 = 7'h5a == _myNewVec_103_T_3[6:0] ? myVec_90 : _GEN_3331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3333 = 7'h5b == _myNewVec_103_T_3[6:0] ? myVec_91 : _GEN_3332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3334 = 7'h5c == _myNewVec_103_T_3[6:0] ? myVec_92 : _GEN_3333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3335 = 7'h5d == _myNewVec_103_T_3[6:0] ? myVec_93 : _GEN_3334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3336 = 7'h5e == _myNewVec_103_T_3[6:0] ? myVec_94 : _GEN_3335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3337 = 7'h5f == _myNewVec_103_T_3[6:0] ? myVec_95 : _GEN_3336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3338 = 7'h60 == _myNewVec_103_T_3[6:0] ? myVec_96 : _GEN_3337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3339 = 7'h61 == _myNewVec_103_T_3[6:0] ? myVec_97 : _GEN_3338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3340 = 7'h62 == _myNewVec_103_T_3[6:0] ? myVec_98 : _GEN_3339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3341 = 7'h63 == _myNewVec_103_T_3[6:0] ? myVec_99 : _GEN_3340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3342 = 7'h64 == _myNewVec_103_T_3[6:0] ? myVec_100 : _GEN_3341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3343 = 7'h65 == _myNewVec_103_T_3[6:0] ? myVec_101 : _GEN_3342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3344 = 7'h66 == _myNewVec_103_T_3[6:0] ? myVec_102 : _GEN_3343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3345 = 7'h67 == _myNewVec_103_T_3[6:0] ? myVec_103 : _GEN_3344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3346 = 7'h68 == _myNewVec_103_T_3[6:0] ? myVec_104 : _GEN_3345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3347 = 7'h69 == _myNewVec_103_T_3[6:0] ? myVec_105 : _GEN_3346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3348 = 7'h6a == _myNewVec_103_T_3[6:0] ? myVec_106 : _GEN_3347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3349 = 7'h6b == _myNewVec_103_T_3[6:0] ? myVec_107 : _GEN_3348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3350 = 7'h6c == _myNewVec_103_T_3[6:0] ? myVec_108 : _GEN_3349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3351 = 7'h6d == _myNewVec_103_T_3[6:0] ? myVec_109 : _GEN_3350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3352 = 7'h6e == _myNewVec_103_T_3[6:0] ? myVec_110 : _GEN_3351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3353 = 7'h6f == _myNewVec_103_T_3[6:0] ? myVec_111 : _GEN_3352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3354 = 7'h70 == _myNewVec_103_T_3[6:0] ? myVec_112 : _GEN_3353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3355 = 7'h71 == _myNewVec_103_T_3[6:0] ? myVec_113 : _GEN_3354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3356 = 7'h72 == _myNewVec_103_T_3[6:0] ? myVec_114 : _GEN_3355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3357 = 7'h73 == _myNewVec_103_T_3[6:0] ? myVec_115 : _GEN_3356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3358 = 7'h74 == _myNewVec_103_T_3[6:0] ? myVec_116 : _GEN_3357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3359 = 7'h75 == _myNewVec_103_T_3[6:0] ? myVec_117 : _GEN_3358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3360 = 7'h76 == _myNewVec_103_T_3[6:0] ? myVec_118 : _GEN_3359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3361 = 7'h77 == _myNewVec_103_T_3[6:0] ? myVec_119 : _GEN_3360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3362 = 7'h78 == _myNewVec_103_T_3[6:0] ? myVec_120 : _GEN_3361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3363 = 7'h79 == _myNewVec_103_T_3[6:0] ? myVec_121 : _GEN_3362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3364 = 7'h7a == _myNewVec_103_T_3[6:0] ? myVec_122 : _GEN_3363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3365 = 7'h7b == _myNewVec_103_T_3[6:0] ? myVec_123 : _GEN_3364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3366 = 7'h7c == _myNewVec_103_T_3[6:0] ? myVec_124 : _GEN_3365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3367 = 7'h7d == _myNewVec_103_T_3[6:0] ? myVec_125 : _GEN_3366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3368 = 7'h7e == _myNewVec_103_T_3[6:0] ? myVec_126 : _GEN_3367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_103 = 7'h7f == _myNewVec_103_T_3[6:0] ? myVec_127 : _GEN_3368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_102_T_3 = _myNewVec_127_T_1 + 16'h19; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3371 = 7'h1 == _myNewVec_102_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3372 = 7'h2 == _myNewVec_102_T_3[6:0] ? myVec_2 : _GEN_3371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3373 = 7'h3 == _myNewVec_102_T_3[6:0] ? myVec_3 : _GEN_3372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3374 = 7'h4 == _myNewVec_102_T_3[6:0] ? myVec_4 : _GEN_3373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3375 = 7'h5 == _myNewVec_102_T_3[6:0] ? myVec_5 : _GEN_3374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3376 = 7'h6 == _myNewVec_102_T_3[6:0] ? myVec_6 : _GEN_3375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3377 = 7'h7 == _myNewVec_102_T_3[6:0] ? myVec_7 : _GEN_3376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3378 = 7'h8 == _myNewVec_102_T_3[6:0] ? myVec_8 : _GEN_3377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3379 = 7'h9 == _myNewVec_102_T_3[6:0] ? myVec_9 : _GEN_3378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3380 = 7'ha == _myNewVec_102_T_3[6:0] ? myVec_10 : _GEN_3379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3381 = 7'hb == _myNewVec_102_T_3[6:0] ? myVec_11 : _GEN_3380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3382 = 7'hc == _myNewVec_102_T_3[6:0] ? myVec_12 : _GEN_3381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3383 = 7'hd == _myNewVec_102_T_3[6:0] ? myVec_13 : _GEN_3382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3384 = 7'he == _myNewVec_102_T_3[6:0] ? myVec_14 : _GEN_3383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3385 = 7'hf == _myNewVec_102_T_3[6:0] ? myVec_15 : _GEN_3384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3386 = 7'h10 == _myNewVec_102_T_3[6:0] ? myVec_16 : _GEN_3385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3387 = 7'h11 == _myNewVec_102_T_3[6:0] ? myVec_17 : _GEN_3386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3388 = 7'h12 == _myNewVec_102_T_3[6:0] ? myVec_18 : _GEN_3387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3389 = 7'h13 == _myNewVec_102_T_3[6:0] ? myVec_19 : _GEN_3388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3390 = 7'h14 == _myNewVec_102_T_3[6:0] ? myVec_20 : _GEN_3389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3391 = 7'h15 == _myNewVec_102_T_3[6:0] ? myVec_21 : _GEN_3390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3392 = 7'h16 == _myNewVec_102_T_3[6:0] ? myVec_22 : _GEN_3391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3393 = 7'h17 == _myNewVec_102_T_3[6:0] ? myVec_23 : _GEN_3392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3394 = 7'h18 == _myNewVec_102_T_3[6:0] ? myVec_24 : _GEN_3393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3395 = 7'h19 == _myNewVec_102_T_3[6:0] ? myVec_25 : _GEN_3394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3396 = 7'h1a == _myNewVec_102_T_3[6:0] ? myVec_26 : _GEN_3395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3397 = 7'h1b == _myNewVec_102_T_3[6:0] ? myVec_27 : _GEN_3396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3398 = 7'h1c == _myNewVec_102_T_3[6:0] ? myVec_28 : _GEN_3397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3399 = 7'h1d == _myNewVec_102_T_3[6:0] ? myVec_29 : _GEN_3398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3400 = 7'h1e == _myNewVec_102_T_3[6:0] ? myVec_30 : _GEN_3399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3401 = 7'h1f == _myNewVec_102_T_3[6:0] ? myVec_31 : _GEN_3400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3402 = 7'h20 == _myNewVec_102_T_3[6:0] ? myVec_32 : _GEN_3401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3403 = 7'h21 == _myNewVec_102_T_3[6:0] ? myVec_33 : _GEN_3402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3404 = 7'h22 == _myNewVec_102_T_3[6:0] ? myVec_34 : _GEN_3403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3405 = 7'h23 == _myNewVec_102_T_3[6:0] ? myVec_35 : _GEN_3404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3406 = 7'h24 == _myNewVec_102_T_3[6:0] ? myVec_36 : _GEN_3405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3407 = 7'h25 == _myNewVec_102_T_3[6:0] ? myVec_37 : _GEN_3406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3408 = 7'h26 == _myNewVec_102_T_3[6:0] ? myVec_38 : _GEN_3407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3409 = 7'h27 == _myNewVec_102_T_3[6:0] ? myVec_39 : _GEN_3408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3410 = 7'h28 == _myNewVec_102_T_3[6:0] ? myVec_40 : _GEN_3409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3411 = 7'h29 == _myNewVec_102_T_3[6:0] ? myVec_41 : _GEN_3410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3412 = 7'h2a == _myNewVec_102_T_3[6:0] ? myVec_42 : _GEN_3411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3413 = 7'h2b == _myNewVec_102_T_3[6:0] ? myVec_43 : _GEN_3412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3414 = 7'h2c == _myNewVec_102_T_3[6:0] ? myVec_44 : _GEN_3413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3415 = 7'h2d == _myNewVec_102_T_3[6:0] ? myVec_45 : _GEN_3414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3416 = 7'h2e == _myNewVec_102_T_3[6:0] ? myVec_46 : _GEN_3415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3417 = 7'h2f == _myNewVec_102_T_3[6:0] ? myVec_47 : _GEN_3416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3418 = 7'h30 == _myNewVec_102_T_3[6:0] ? myVec_48 : _GEN_3417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3419 = 7'h31 == _myNewVec_102_T_3[6:0] ? myVec_49 : _GEN_3418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3420 = 7'h32 == _myNewVec_102_T_3[6:0] ? myVec_50 : _GEN_3419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3421 = 7'h33 == _myNewVec_102_T_3[6:0] ? myVec_51 : _GEN_3420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3422 = 7'h34 == _myNewVec_102_T_3[6:0] ? myVec_52 : _GEN_3421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3423 = 7'h35 == _myNewVec_102_T_3[6:0] ? myVec_53 : _GEN_3422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3424 = 7'h36 == _myNewVec_102_T_3[6:0] ? myVec_54 : _GEN_3423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3425 = 7'h37 == _myNewVec_102_T_3[6:0] ? myVec_55 : _GEN_3424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3426 = 7'h38 == _myNewVec_102_T_3[6:0] ? myVec_56 : _GEN_3425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3427 = 7'h39 == _myNewVec_102_T_3[6:0] ? myVec_57 : _GEN_3426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3428 = 7'h3a == _myNewVec_102_T_3[6:0] ? myVec_58 : _GEN_3427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3429 = 7'h3b == _myNewVec_102_T_3[6:0] ? myVec_59 : _GEN_3428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3430 = 7'h3c == _myNewVec_102_T_3[6:0] ? myVec_60 : _GEN_3429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3431 = 7'h3d == _myNewVec_102_T_3[6:0] ? myVec_61 : _GEN_3430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3432 = 7'h3e == _myNewVec_102_T_3[6:0] ? myVec_62 : _GEN_3431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3433 = 7'h3f == _myNewVec_102_T_3[6:0] ? myVec_63 : _GEN_3432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3434 = 7'h40 == _myNewVec_102_T_3[6:0] ? myVec_64 : _GEN_3433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3435 = 7'h41 == _myNewVec_102_T_3[6:0] ? myVec_65 : _GEN_3434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3436 = 7'h42 == _myNewVec_102_T_3[6:0] ? myVec_66 : _GEN_3435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3437 = 7'h43 == _myNewVec_102_T_3[6:0] ? myVec_67 : _GEN_3436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3438 = 7'h44 == _myNewVec_102_T_3[6:0] ? myVec_68 : _GEN_3437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3439 = 7'h45 == _myNewVec_102_T_3[6:0] ? myVec_69 : _GEN_3438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3440 = 7'h46 == _myNewVec_102_T_3[6:0] ? myVec_70 : _GEN_3439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3441 = 7'h47 == _myNewVec_102_T_3[6:0] ? myVec_71 : _GEN_3440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3442 = 7'h48 == _myNewVec_102_T_3[6:0] ? myVec_72 : _GEN_3441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3443 = 7'h49 == _myNewVec_102_T_3[6:0] ? myVec_73 : _GEN_3442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3444 = 7'h4a == _myNewVec_102_T_3[6:0] ? myVec_74 : _GEN_3443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3445 = 7'h4b == _myNewVec_102_T_3[6:0] ? myVec_75 : _GEN_3444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3446 = 7'h4c == _myNewVec_102_T_3[6:0] ? myVec_76 : _GEN_3445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3447 = 7'h4d == _myNewVec_102_T_3[6:0] ? myVec_77 : _GEN_3446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3448 = 7'h4e == _myNewVec_102_T_3[6:0] ? myVec_78 : _GEN_3447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3449 = 7'h4f == _myNewVec_102_T_3[6:0] ? myVec_79 : _GEN_3448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3450 = 7'h50 == _myNewVec_102_T_3[6:0] ? myVec_80 : _GEN_3449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3451 = 7'h51 == _myNewVec_102_T_3[6:0] ? myVec_81 : _GEN_3450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3452 = 7'h52 == _myNewVec_102_T_3[6:0] ? myVec_82 : _GEN_3451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3453 = 7'h53 == _myNewVec_102_T_3[6:0] ? myVec_83 : _GEN_3452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3454 = 7'h54 == _myNewVec_102_T_3[6:0] ? myVec_84 : _GEN_3453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3455 = 7'h55 == _myNewVec_102_T_3[6:0] ? myVec_85 : _GEN_3454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3456 = 7'h56 == _myNewVec_102_T_3[6:0] ? myVec_86 : _GEN_3455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3457 = 7'h57 == _myNewVec_102_T_3[6:0] ? myVec_87 : _GEN_3456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3458 = 7'h58 == _myNewVec_102_T_3[6:0] ? myVec_88 : _GEN_3457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3459 = 7'h59 == _myNewVec_102_T_3[6:0] ? myVec_89 : _GEN_3458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3460 = 7'h5a == _myNewVec_102_T_3[6:0] ? myVec_90 : _GEN_3459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3461 = 7'h5b == _myNewVec_102_T_3[6:0] ? myVec_91 : _GEN_3460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3462 = 7'h5c == _myNewVec_102_T_3[6:0] ? myVec_92 : _GEN_3461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3463 = 7'h5d == _myNewVec_102_T_3[6:0] ? myVec_93 : _GEN_3462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3464 = 7'h5e == _myNewVec_102_T_3[6:0] ? myVec_94 : _GEN_3463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3465 = 7'h5f == _myNewVec_102_T_3[6:0] ? myVec_95 : _GEN_3464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3466 = 7'h60 == _myNewVec_102_T_3[6:0] ? myVec_96 : _GEN_3465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3467 = 7'h61 == _myNewVec_102_T_3[6:0] ? myVec_97 : _GEN_3466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3468 = 7'h62 == _myNewVec_102_T_3[6:0] ? myVec_98 : _GEN_3467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3469 = 7'h63 == _myNewVec_102_T_3[6:0] ? myVec_99 : _GEN_3468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3470 = 7'h64 == _myNewVec_102_T_3[6:0] ? myVec_100 : _GEN_3469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3471 = 7'h65 == _myNewVec_102_T_3[6:0] ? myVec_101 : _GEN_3470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3472 = 7'h66 == _myNewVec_102_T_3[6:0] ? myVec_102 : _GEN_3471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3473 = 7'h67 == _myNewVec_102_T_3[6:0] ? myVec_103 : _GEN_3472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3474 = 7'h68 == _myNewVec_102_T_3[6:0] ? myVec_104 : _GEN_3473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3475 = 7'h69 == _myNewVec_102_T_3[6:0] ? myVec_105 : _GEN_3474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3476 = 7'h6a == _myNewVec_102_T_3[6:0] ? myVec_106 : _GEN_3475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3477 = 7'h6b == _myNewVec_102_T_3[6:0] ? myVec_107 : _GEN_3476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3478 = 7'h6c == _myNewVec_102_T_3[6:0] ? myVec_108 : _GEN_3477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3479 = 7'h6d == _myNewVec_102_T_3[6:0] ? myVec_109 : _GEN_3478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3480 = 7'h6e == _myNewVec_102_T_3[6:0] ? myVec_110 : _GEN_3479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3481 = 7'h6f == _myNewVec_102_T_3[6:0] ? myVec_111 : _GEN_3480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3482 = 7'h70 == _myNewVec_102_T_3[6:0] ? myVec_112 : _GEN_3481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3483 = 7'h71 == _myNewVec_102_T_3[6:0] ? myVec_113 : _GEN_3482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3484 = 7'h72 == _myNewVec_102_T_3[6:0] ? myVec_114 : _GEN_3483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3485 = 7'h73 == _myNewVec_102_T_3[6:0] ? myVec_115 : _GEN_3484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3486 = 7'h74 == _myNewVec_102_T_3[6:0] ? myVec_116 : _GEN_3485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3487 = 7'h75 == _myNewVec_102_T_3[6:0] ? myVec_117 : _GEN_3486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3488 = 7'h76 == _myNewVec_102_T_3[6:0] ? myVec_118 : _GEN_3487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3489 = 7'h77 == _myNewVec_102_T_3[6:0] ? myVec_119 : _GEN_3488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3490 = 7'h78 == _myNewVec_102_T_3[6:0] ? myVec_120 : _GEN_3489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3491 = 7'h79 == _myNewVec_102_T_3[6:0] ? myVec_121 : _GEN_3490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3492 = 7'h7a == _myNewVec_102_T_3[6:0] ? myVec_122 : _GEN_3491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3493 = 7'h7b == _myNewVec_102_T_3[6:0] ? myVec_123 : _GEN_3492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3494 = 7'h7c == _myNewVec_102_T_3[6:0] ? myVec_124 : _GEN_3493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3495 = 7'h7d == _myNewVec_102_T_3[6:0] ? myVec_125 : _GEN_3494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3496 = 7'h7e == _myNewVec_102_T_3[6:0] ? myVec_126 : _GEN_3495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_102 = 7'h7f == _myNewVec_102_T_3[6:0] ? myVec_127 : _GEN_3496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_101_T_3 = _myNewVec_127_T_1 + 16'h1a; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3499 = 7'h1 == _myNewVec_101_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3500 = 7'h2 == _myNewVec_101_T_3[6:0] ? myVec_2 : _GEN_3499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3501 = 7'h3 == _myNewVec_101_T_3[6:0] ? myVec_3 : _GEN_3500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3502 = 7'h4 == _myNewVec_101_T_3[6:0] ? myVec_4 : _GEN_3501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3503 = 7'h5 == _myNewVec_101_T_3[6:0] ? myVec_5 : _GEN_3502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3504 = 7'h6 == _myNewVec_101_T_3[6:0] ? myVec_6 : _GEN_3503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3505 = 7'h7 == _myNewVec_101_T_3[6:0] ? myVec_7 : _GEN_3504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3506 = 7'h8 == _myNewVec_101_T_3[6:0] ? myVec_8 : _GEN_3505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3507 = 7'h9 == _myNewVec_101_T_3[6:0] ? myVec_9 : _GEN_3506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3508 = 7'ha == _myNewVec_101_T_3[6:0] ? myVec_10 : _GEN_3507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3509 = 7'hb == _myNewVec_101_T_3[6:0] ? myVec_11 : _GEN_3508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3510 = 7'hc == _myNewVec_101_T_3[6:0] ? myVec_12 : _GEN_3509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3511 = 7'hd == _myNewVec_101_T_3[6:0] ? myVec_13 : _GEN_3510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3512 = 7'he == _myNewVec_101_T_3[6:0] ? myVec_14 : _GEN_3511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3513 = 7'hf == _myNewVec_101_T_3[6:0] ? myVec_15 : _GEN_3512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3514 = 7'h10 == _myNewVec_101_T_3[6:0] ? myVec_16 : _GEN_3513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3515 = 7'h11 == _myNewVec_101_T_3[6:0] ? myVec_17 : _GEN_3514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3516 = 7'h12 == _myNewVec_101_T_3[6:0] ? myVec_18 : _GEN_3515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3517 = 7'h13 == _myNewVec_101_T_3[6:0] ? myVec_19 : _GEN_3516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3518 = 7'h14 == _myNewVec_101_T_3[6:0] ? myVec_20 : _GEN_3517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3519 = 7'h15 == _myNewVec_101_T_3[6:0] ? myVec_21 : _GEN_3518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3520 = 7'h16 == _myNewVec_101_T_3[6:0] ? myVec_22 : _GEN_3519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3521 = 7'h17 == _myNewVec_101_T_3[6:0] ? myVec_23 : _GEN_3520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3522 = 7'h18 == _myNewVec_101_T_3[6:0] ? myVec_24 : _GEN_3521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3523 = 7'h19 == _myNewVec_101_T_3[6:0] ? myVec_25 : _GEN_3522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3524 = 7'h1a == _myNewVec_101_T_3[6:0] ? myVec_26 : _GEN_3523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3525 = 7'h1b == _myNewVec_101_T_3[6:0] ? myVec_27 : _GEN_3524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3526 = 7'h1c == _myNewVec_101_T_3[6:0] ? myVec_28 : _GEN_3525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3527 = 7'h1d == _myNewVec_101_T_3[6:0] ? myVec_29 : _GEN_3526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3528 = 7'h1e == _myNewVec_101_T_3[6:0] ? myVec_30 : _GEN_3527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3529 = 7'h1f == _myNewVec_101_T_3[6:0] ? myVec_31 : _GEN_3528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3530 = 7'h20 == _myNewVec_101_T_3[6:0] ? myVec_32 : _GEN_3529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3531 = 7'h21 == _myNewVec_101_T_3[6:0] ? myVec_33 : _GEN_3530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3532 = 7'h22 == _myNewVec_101_T_3[6:0] ? myVec_34 : _GEN_3531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3533 = 7'h23 == _myNewVec_101_T_3[6:0] ? myVec_35 : _GEN_3532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3534 = 7'h24 == _myNewVec_101_T_3[6:0] ? myVec_36 : _GEN_3533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3535 = 7'h25 == _myNewVec_101_T_3[6:0] ? myVec_37 : _GEN_3534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3536 = 7'h26 == _myNewVec_101_T_3[6:0] ? myVec_38 : _GEN_3535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3537 = 7'h27 == _myNewVec_101_T_3[6:0] ? myVec_39 : _GEN_3536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3538 = 7'h28 == _myNewVec_101_T_3[6:0] ? myVec_40 : _GEN_3537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3539 = 7'h29 == _myNewVec_101_T_3[6:0] ? myVec_41 : _GEN_3538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3540 = 7'h2a == _myNewVec_101_T_3[6:0] ? myVec_42 : _GEN_3539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3541 = 7'h2b == _myNewVec_101_T_3[6:0] ? myVec_43 : _GEN_3540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3542 = 7'h2c == _myNewVec_101_T_3[6:0] ? myVec_44 : _GEN_3541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3543 = 7'h2d == _myNewVec_101_T_3[6:0] ? myVec_45 : _GEN_3542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3544 = 7'h2e == _myNewVec_101_T_3[6:0] ? myVec_46 : _GEN_3543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3545 = 7'h2f == _myNewVec_101_T_3[6:0] ? myVec_47 : _GEN_3544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3546 = 7'h30 == _myNewVec_101_T_3[6:0] ? myVec_48 : _GEN_3545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3547 = 7'h31 == _myNewVec_101_T_3[6:0] ? myVec_49 : _GEN_3546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3548 = 7'h32 == _myNewVec_101_T_3[6:0] ? myVec_50 : _GEN_3547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3549 = 7'h33 == _myNewVec_101_T_3[6:0] ? myVec_51 : _GEN_3548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3550 = 7'h34 == _myNewVec_101_T_3[6:0] ? myVec_52 : _GEN_3549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3551 = 7'h35 == _myNewVec_101_T_3[6:0] ? myVec_53 : _GEN_3550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3552 = 7'h36 == _myNewVec_101_T_3[6:0] ? myVec_54 : _GEN_3551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3553 = 7'h37 == _myNewVec_101_T_3[6:0] ? myVec_55 : _GEN_3552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3554 = 7'h38 == _myNewVec_101_T_3[6:0] ? myVec_56 : _GEN_3553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3555 = 7'h39 == _myNewVec_101_T_3[6:0] ? myVec_57 : _GEN_3554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3556 = 7'h3a == _myNewVec_101_T_3[6:0] ? myVec_58 : _GEN_3555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3557 = 7'h3b == _myNewVec_101_T_3[6:0] ? myVec_59 : _GEN_3556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3558 = 7'h3c == _myNewVec_101_T_3[6:0] ? myVec_60 : _GEN_3557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3559 = 7'h3d == _myNewVec_101_T_3[6:0] ? myVec_61 : _GEN_3558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3560 = 7'h3e == _myNewVec_101_T_3[6:0] ? myVec_62 : _GEN_3559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3561 = 7'h3f == _myNewVec_101_T_3[6:0] ? myVec_63 : _GEN_3560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3562 = 7'h40 == _myNewVec_101_T_3[6:0] ? myVec_64 : _GEN_3561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3563 = 7'h41 == _myNewVec_101_T_3[6:0] ? myVec_65 : _GEN_3562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3564 = 7'h42 == _myNewVec_101_T_3[6:0] ? myVec_66 : _GEN_3563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3565 = 7'h43 == _myNewVec_101_T_3[6:0] ? myVec_67 : _GEN_3564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3566 = 7'h44 == _myNewVec_101_T_3[6:0] ? myVec_68 : _GEN_3565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3567 = 7'h45 == _myNewVec_101_T_3[6:0] ? myVec_69 : _GEN_3566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3568 = 7'h46 == _myNewVec_101_T_3[6:0] ? myVec_70 : _GEN_3567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3569 = 7'h47 == _myNewVec_101_T_3[6:0] ? myVec_71 : _GEN_3568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3570 = 7'h48 == _myNewVec_101_T_3[6:0] ? myVec_72 : _GEN_3569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3571 = 7'h49 == _myNewVec_101_T_3[6:0] ? myVec_73 : _GEN_3570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3572 = 7'h4a == _myNewVec_101_T_3[6:0] ? myVec_74 : _GEN_3571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3573 = 7'h4b == _myNewVec_101_T_3[6:0] ? myVec_75 : _GEN_3572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3574 = 7'h4c == _myNewVec_101_T_3[6:0] ? myVec_76 : _GEN_3573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3575 = 7'h4d == _myNewVec_101_T_3[6:0] ? myVec_77 : _GEN_3574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3576 = 7'h4e == _myNewVec_101_T_3[6:0] ? myVec_78 : _GEN_3575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3577 = 7'h4f == _myNewVec_101_T_3[6:0] ? myVec_79 : _GEN_3576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3578 = 7'h50 == _myNewVec_101_T_3[6:0] ? myVec_80 : _GEN_3577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3579 = 7'h51 == _myNewVec_101_T_3[6:0] ? myVec_81 : _GEN_3578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3580 = 7'h52 == _myNewVec_101_T_3[6:0] ? myVec_82 : _GEN_3579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3581 = 7'h53 == _myNewVec_101_T_3[6:0] ? myVec_83 : _GEN_3580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3582 = 7'h54 == _myNewVec_101_T_3[6:0] ? myVec_84 : _GEN_3581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3583 = 7'h55 == _myNewVec_101_T_3[6:0] ? myVec_85 : _GEN_3582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3584 = 7'h56 == _myNewVec_101_T_3[6:0] ? myVec_86 : _GEN_3583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3585 = 7'h57 == _myNewVec_101_T_3[6:0] ? myVec_87 : _GEN_3584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3586 = 7'h58 == _myNewVec_101_T_3[6:0] ? myVec_88 : _GEN_3585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3587 = 7'h59 == _myNewVec_101_T_3[6:0] ? myVec_89 : _GEN_3586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3588 = 7'h5a == _myNewVec_101_T_3[6:0] ? myVec_90 : _GEN_3587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3589 = 7'h5b == _myNewVec_101_T_3[6:0] ? myVec_91 : _GEN_3588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3590 = 7'h5c == _myNewVec_101_T_3[6:0] ? myVec_92 : _GEN_3589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3591 = 7'h5d == _myNewVec_101_T_3[6:0] ? myVec_93 : _GEN_3590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3592 = 7'h5e == _myNewVec_101_T_3[6:0] ? myVec_94 : _GEN_3591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3593 = 7'h5f == _myNewVec_101_T_3[6:0] ? myVec_95 : _GEN_3592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3594 = 7'h60 == _myNewVec_101_T_3[6:0] ? myVec_96 : _GEN_3593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3595 = 7'h61 == _myNewVec_101_T_3[6:0] ? myVec_97 : _GEN_3594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3596 = 7'h62 == _myNewVec_101_T_3[6:0] ? myVec_98 : _GEN_3595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3597 = 7'h63 == _myNewVec_101_T_3[6:0] ? myVec_99 : _GEN_3596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3598 = 7'h64 == _myNewVec_101_T_3[6:0] ? myVec_100 : _GEN_3597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3599 = 7'h65 == _myNewVec_101_T_3[6:0] ? myVec_101 : _GEN_3598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3600 = 7'h66 == _myNewVec_101_T_3[6:0] ? myVec_102 : _GEN_3599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3601 = 7'h67 == _myNewVec_101_T_3[6:0] ? myVec_103 : _GEN_3600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3602 = 7'h68 == _myNewVec_101_T_3[6:0] ? myVec_104 : _GEN_3601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3603 = 7'h69 == _myNewVec_101_T_3[6:0] ? myVec_105 : _GEN_3602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3604 = 7'h6a == _myNewVec_101_T_3[6:0] ? myVec_106 : _GEN_3603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3605 = 7'h6b == _myNewVec_101_T_3[6:0] ? myVec_107 : _GEN_3604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3606 = 7'h6c == _myNewVec_101_T_3[6:0] ? myVec_108 : _GEN_3605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3607 = 7'h6d == _myNewVec_101_T_3[6:0] ? myVec_109 : _GEN_3606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3608 = 7'h6e == _myNewVec_101_T_3[6:0] ? myVec_110 : _GEN_3607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3609 = 7'h6f == _myNewVec_101_T_3[6:0] ? myVec_111 : _GEN_3608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3610 = 7'h70 == _myNewVec_101_T_3[6:0] ? myVec_112 : _GEN_3609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3611 = 7'h71 == _myNewVec_101_T_3[6:0] ? myVec_113 : _GEN_3610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3612 = 7'h72 == _myNewVec_101_T_3[6:0] ? myVec_114 : _GEN_3611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3613 = 7'h73 == _myNewVec_101_T_3[6:0] ? myVec_115 : _GEN_3612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3614 = 7'h74 == _myNewVec_101_T_3[6:0] ? myVec_116 : _GEN_3613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3615 = 7'h75 == _myNewVec_101_T_3[6:0] ? myVec_117 : _GEN_3614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3616 = 7'h76 == _myNewVec_101_T_3[6:0] ? myVec_118 : _GEN_3615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3617 = 7'h77 == _myNewVec_101_T_3[6:0] ? myVec_119 : _GEN_3616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3618 = 7'h78 == _myNewVec_101_T_3[6:0] ? myVec_120 : _GEN_3617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3619 = 7'h79 == _myNewVec_101_T_3[6:0] ? myVec_121 : _GEN_3618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3620 = 7'h7a == _myNewVec_101_T_3[6:0] ? myVec_122 : _GEN_3619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3621 = 7'h7b == _myNewVec_101_T_3[6:0] ? myVec_123 : _GEN_3620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3622 = 7'h7c == _myNewVec_101_T_3[6:0] ? myVec_124 : _GEN_3621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3623 = 7'h7d == _myNewVec_101_T_3[6:0] ? myVec_125 : _GEN_3622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3624 = 7'h7e == _myNewVec_101_T_3[6:0] ? myVec_126 : _GEN_3623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_101 = 7'h7f == _myNewVec_101_T_3[6:0] ? myVec_127 : _GEN_3624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_100_T_3 = _myNewVec_127_T_1 + 16'h1b; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3627 = 7'h1 == _myNewVec_100_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3628 = 7'h2 == _myNewVec_100_T_3[6:0] ? myVec_2 : _GEN_3627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3629 = 7'h3 == _myNewVec_100_T_3[6:0] ? myVec_3 : _GEN_3628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3630 = 7'h4 == _myNewVec_100_T_3[6:0] ? myVec_4 : _GEN_3629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3631 = 7'h5 == _myNewVec_100_T_3[6:0] ? myVec_5 : _GEN_3630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3632 = 7'h6 == _myNewVec_100_T_3[6:0] ? myVec_6 : _GEN_3631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3633 = 7'h7 == _myNewVec_100_T_3[6:0] ? myVec_7 : _GEN_3632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3634 = 7'h8 == _myNewVec_100_T_3[6:0] ? myVec_8 : _GEN_3633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3635 = 7'h9 == _myNewVec_100_T_3[6:0] ? myVec_9 : _GEN_3634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3636 = 7'ha == _myNewVec_100_T_3[6:0] ? myVec_10 : _GEN_3635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3637 = 7'hb == _myNewVec_100_T_3[6:0] ? myVec_11 : _GEN_3636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3638 = 7'hc == _myNewVec_100_T_3[6:0] ? myVec_12 : _GEN_3637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3639 = 7'hd == _myNewVec_100_T_3[6:0] ? myVec_13 : _GEN_3638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3640 = 7'he == _myNewVec_100_T_3[6:0] ? myVec_14 : _GEN_3639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3641 = 7'hf == _myNewVec_100_T_3[6:0] ? myVec_15 : _GEN_3640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3642 = 7'h10 == _myNewVec_100_T_3[6:0] ? myVec_16 : _GEN_3641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3643 = 7'h11 == _myNewVec_100_T_3[6:0] ? myVec_17 : _GEN_3642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3644 = 7'h12 == _myNewVec_100_T_3[6:0] ? myVec_18 : _GEN_3643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3645 = 7'h13 == _myNewVec_100_T_3[6:0] ? myVec_19 : _GEN_3644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3646 = 7'h14 == _myNewVec_100_T_3[6:0] ? myVec_20 : _GEN_3645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3647 = 7'h15 == _myNewVec_100_T_3[6:0] ? myVec_21 : _GEN_3646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3648 = 7'h16 == _myNewVec_100_T_3[6:0] ? myVec_22 : _GEN_3647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3649 = 7'h17 == _myNewVec_100_T_3[6:0] ? myVec_23 : _GEN_3648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3650 = 7'h18 == _myNewVec_100_T_3[6:0] ? myVec_24 : _GEN_3649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3651 = 7'h19 == _myNewVec_100_T_3[6:0] ? myVec_25 : _GEN_3650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3652 = 7'h1a == _myNewVec_100_T_3[6:0] ? myVec_26 : _GEN_3651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3653 = 7'h1b == _myNewVec_100_T_3[6:0] ? myVec_27 : _GEN_3652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3654 = 7'h1c == _myNewVec_100_T_3[6:0] ? myVec_28 : _GEN_3653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3655 = 7'h1d == _myNewVec_100_T_3[6:0] ? myVec_29 : _GEN_3654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3656 = 7'h1e == _myNewVec_100_T_3[6:0] ? myVec_30 : _GEN_3655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3657 = 7'h1f == _myNewVec_100_T_3[6:0] ? myVec_31 : _GEN_3656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3658 = 7'h20 == _myNewVec_100_T_3[6:0] ? myVec_32 : _GEN_3657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3659 = 7'h21 == _myNewVec_100_T_3[6:0] ? myVec_33 : _GEN_3658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3660 = 7'h22 == _myNewVec_100_T_3[6:0] ? myVec_34 : _GEN_3659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3661 = 7'h23 == _myNewVec_100_T_3[6:0] ? myVec_35 : _GEN_3660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3662 = 7'h24 == _myNewVec_100_T_3[6:0] ? myVec_36 : _GEN_3661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3663 = 7'h25 == _myNewVec_100_T_3[6:0] ? myVec_37 : _GEN_3662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3664 = 7'h26 == _myNewVec_100_T_3[6:0] ? myVec_38 : _GEN_3663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3665 = 7'h27 == _myNewVec_100_T_3[6:0] ? myVec_39 : _GEN_3664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3666 = 7'h28 == _myNewVec_100_T_3[6:0] ? myVec_40 : _GEN_3665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3667 = 7'h29 == _myNewVec_100_T_3[6:0] ? myVec_41 : _GEN_3666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3668 = 7'h2a == _myNewVec_100_T_3[6:0] ? myVec_42 : _GEN_3667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3669 = 7'h2b == _myNewVec_100_T_3[6:0] ? myVec_43 : _GEN_3668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3670 = 7'h2c == _myNewVec_100_T_3[6:0] ? myVec_44 : _GEN_3669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3671 = 7'h2d == _myNewVec_100_T_3[6:0] ? myVec_45 : _GEN_3670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3672 = 7'h2e == _myNewVec_100_T_3[6:0] ? myVec_46 : _GEN_3671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3673 = 7'h2f == _myNewVec_100_T_3[6:0] ? myVec_47 : _GEN_3672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3674 = 7'h30 == _myNewVec_100_T_3[6:0] ? myVec_48 : _GEN_3673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3675 = 7'h31 == _myNewVec_100_T_3[6:0] ? myVec_49 : _GEN_3674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3676 = 7'h32 == _myNewVec_100_T_3[6:0] ? myVec_50 : _GEN_3675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3677 = 7'h33 == _myNewVec_100_T_3[6:0] ? myVec_51 : _GEN_3676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3678 = 7'h34 == _myNewVec_100_T_3[6:0] ? myVec_52 : _GEN_3677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3679 = 7'h35 == _myNewVec_100_T_3[6:0] ? myVec_53 : _GEN_3678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3680 = 7'h36 == _myNewVec_100_T_3[6:0] ? myVec_54 : _GEN_3679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3681 = 7'h37 == _myNewVec_100_T_3[6:0] ? myVec_55 : _GEN_3680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3682 = 7'h38 == _myNewVec_100_T_3[6:0] ? myVec_56 : _GEN_3681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3683 = 7'h39 == _myNewVec_100_T_3[6:0] ? myVec_57 : _GEN_3682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3684 = 7'h3a == _myNewVec_100_T_3[6:0] ? myVec_58 : _GEN_3683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3685 = 7'h3b == _myNewVec_100_T_3[6:0] ? myVec_59 : _GEN_3684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3686 = 7'h3c == _myNewVec_100_T_3[6:0] ? myVec_60 : _GEN_3685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3687 = 7'h3d == _myNewVec_100_T_3[6:0] ? myVec_61 : _GEN_3686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3688 = 7'h3e == _myNewVec_100_T_3[6:0] ? myVec_62 : _GEN_3687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3689 = 7'h3f == _myNewVec_100_T_3[6:0] ? myVec_63 : _GEN_3688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3690 = 7'h40 == _myNewVec_100_T_3[6:0] ? myVec_64 : _GEN_3689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3691 = 7'h41 == _myNewVec_100_T_3[6:0] ? myVec_65 : _GEN_3690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3692 = 7'h42 == _myNewVec_100_T_3[6:0] ? myVec_66 : _GEN_3691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3693 = 7'h43 == _myNewVec_100_T_3[6:0] ? myVec_67 : _GEN_3692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3694 = 7'h44 == _myNewVec_100_T_3[6:0] ? myVec_68 : _GEN_3693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3695 = 7'h45 == _myNewVec_100_T_3[6:0] ? myVec_69 : _GEN_3694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3696 = 7'h46 == _myNewVec_100_T_3[6:0] ? myVec_70 : _GEN_3695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3697 = 7'h47 == _myNewVec_100_T_3[6:0] ? myVec_71 : _GEN_3696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3698 = 7'h48 == _myNewVec_100_T_3[6:0] ? myVec_72 : _GEN_3697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3699 = 7'h49 == _myNewVec_100_T_3[6:0] ? myVec_73 : _GEN_3698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3700 = 7'h4a == _myNewVec_100_T_3[6:0] ? myVec_74 : _GEN_3699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3701 = 7'h4b == _myNewVec_100_T_3[6:0] ? myVec_75 : _GEN_3700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3702 = 7'h4c == _myNewVec_100_T_3[6:0] ? myVec_76 : _GEN_3701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3703 = 7'h4d == _myNewVec_100_T_3[6:0] ? myVec_77 : _GEN_3702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3704 = 7'h4e == _myNewVec_100_T_3[6:0] ? myVec_78 : _GEN_3703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3705 = 7'h4f == _myNewVec_100_T_3[6:0] ? myVec_79 : _GEN_3704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3706 = 7'h50 == _myNewVec_100_T_3[6:0] ? myVec_80 : _GEN_3705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3707 = 7'h51 == _myNewVec_100_T_3[6:0] ? myVec_81 : _GEN_3706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3708 = 7'h52 == _myNewVec_100_T_3[6:0] ? myVec_82 : _GEN_3707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3709 = 7'h53 == _myNewVec_100_T_3[6:0] ? myVec_83 : _GEN_3708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3710 = 7'h54 == _myNewVec_100_T_3[6:0] ? myVec_84 : _GEN_3709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3711 = 7'h55 == _myNewVec_100_T_3[6:0] ? myVec_85 : _GEN_3710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3712 = 7'h56 == _myNewVec_100_T_3[6:0] ? myVec_86 : _GEN_3711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3713 = 7'h57 == _myNewVec_100_T_3[6:0] ? myVec_87 : _GEN_3712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3714 = 7'h58 == _myNewVec_100_T_3[6:0] ? myVec_88 : _GEN_3713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3715 = 7'h59 == _myNewVec_100_T_3[6:0] ? myVec_89 : _GEN_3714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3716 = 7'h5a == _myNewVec_100_T_3[6:0] ? myVec_90 : _GEN_3715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3717 = 7'h5b == _myNewVec_100_T_3[6:0] ? myVec_91 : _GEN_3716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3718 = 7'h5c == _myNewVec_100_T_3[6:0] ? myVec_92 : _GEN_3717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3719 = 7'h5d == _myNewVec_100_T_3[6:0] ? myVec_93 : _GEN_3718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3720 = 7'h5e == _myNewVec_100_T_3[6:0] ? myVec_94 : _GEN_3719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3721 = 7'h5f == _myNewVec_100_T_3[6:0] ? myVec_95 : _GEN_3720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3722 = 7'h60 == _myNewVec_100_T_3[6:0] ? myVec_96 : _GEN_3721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3723 = 7'h61 == _myNewVec_100_T_3[6:0] ? myVec_97 : _GEN_3722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3724 = 7'h62 == _myNewVec_100_T_3[6:0] ? myVec_98 : _GEN_3723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3725 = 7'h63 == _myNewVec_100_T_3[6:0] ? myVec_99 : _GEN_3724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3726 = 7'h64 == _myNewVec_100_T_3[6:0] ? myVec_100 : _GEN_3725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3727 = 7'h65 == _myNewVec_100_T_3[6:0] ? myVec_101 : _GEN_3726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3728 = 7'h66 == _myNewVec_100_T_3[6:0] ? myVec_102 : _GEN_3727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3729 = 7'h67 == _myNewVec_100_T_3[6:0] ? myVec_103 : _GEN_3728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3730 = 7'h68 == _myNewVec_100_T_3[6:0] ? myVec_104 : _GEN_3729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3731 = 7'h69 == _myNewVec_100_T_3[6:0] ? myVec_105 : _GEN_3730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3732 = 7'h6a == _myNewVec_100_T_3[6:0] ? myVec_106 : _GEN_3731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3733 = 7'h6b == _myNewVec_100_T_3[6:0] ? myVec_107 : _GEN_3732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3734 = 7'h6c == _myNewVec_100_T_3[6:0] ? myVec_108 : _GEN_3733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3735 = 7'h6d == _myNewVec_100_T_3[6:0] ? myVec_109 : _GEN_3734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3736 = 7'h6e == _myNewVec_100_T_3[6:0] ? myVec_110 : _GEN_3735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3737 = 7'h6f == _myNewVec_100_T_3[6:0] ? myVec_111 : _GEN_3736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3738 = 7'h70 == _myNewVec_100_T_3[6:0] ? myVec_112 : _GEN_3737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3739 = 7'h71 == _myNewVec_100_T_3[6:0] ? myVec_113 : _GEN_3738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3740 = 7'h72 == _myNewVec_100_T_3[6:0] ? myVec_114 : _GEN_3739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3741 = 7'h73 == _myNewVec_100_T_3[6:0] ? myVec_115 : _GEN_3740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3742 = 7'h74 == _myNewVec_100_T_3[6:0] ? myVec_116 : _GEN_3741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3743 = 7'h75 == _myNewVec_100_T_3[6:0] ? myVec_117 : _GEN_3742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3744 = 7'h76 == _myNewVec_100_T_3[6:0] ? myVec_118 : _GEN_3743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3745 = 7'h77 == _myNewVec_100_T_3[6:0] ? myVec_119 : _GEN_3744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3746 = 7'h78 == _myNewVec_100_T_3[6:0] ? myVec_120 : _GEN_3745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3747 = 7'h79 == _myNewVec_100_T_3[6:0] ? myVec_121 : _GEN_3746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3748 = 7'h7a == _myNewVec_100_T_3[6:0] ? myVec_122 : _GEN_3747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3749 = 7'h7b == _myNewVec_100_T_3[6:0] ? myVec_123 : _GEN_3748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3750 = 7'h7c == _myNewVec_100_T_3[6:0] ? myVec_124 : _GEN_3749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3751 = 7'h7d == _myNewVec_100_T_3[6:0] ? myVec_125 : _GEN_3750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3752 = 7'h7e == _myNewVec_100_T_3[6:0] ? myVec_126 : _GEN_3751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_100 = 7'h7f == _myNewVec_100_T_3[6:0] ? myVec_127 : _GEN_3752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_99_T_3 = _myNewVec_127_T_1 + 16'h1c; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3755 = 7'h1 == _myNewVec_99_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3756 = 7'h2 == _myNewVec_99_T_3[6:0] ? myVec_2 : _GEN_3755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3757 = 7'h3 == _myNewVec_99_T_3[6:0] ? myVec_3 : _GEN_3756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3758 = 7'h4 == _myNewVec_99_T_3[6:0] ? myVec_4 : _GEN_3757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3759 = 7'h5 == _myNewVec_99_T_3[6:0] ? myVec_5 : _GEN_3758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3760 = 7'h6 == _myNewVec_99_T_3[6:0] ? myVec_6 : _GEN_3759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3761 = 7'h7 == _myNewVec_99_T_3[6:0] ? myVec_7 : _GEN_3760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3762 = 7'h8 == _myNewVec_99_T_3[6:0] ? myVec_8 : _GEN_3761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3763 = 7'h9 == _myNewVec_99_T_3[6:0] ? myVec_9 : _GEN_3762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3764 = 7'ha == _myNewVec_99_T_3[6:0] ? myVec_10 : _GEN_3763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3765 = 7'hb == _myNewVec_99_T_3[6:0] ? myVec_11 : _GEN_3764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3766 = 7'hc == _myNewVec_99_T_3[6:0] ? myVec_12 : _GEN_3765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3767 = 7'hd == _myNewVec_99_T_3[6:0] ? myVec_13 : _GEN_3766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3768 = 7'he == _myNewVec_99_T_3[6:0] ? myVec_14 : _GEN_3767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3769 = 7'hf == _myNewVec_99_T_3[6:0] ? myVec_15 : _GEN_3768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3770 = 7'h10 == _myNewVec_99_T_3[6:0] ? myVec_16 : _GEN_3769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3771 = 7'h11 == _myNewVec_99_T_3[6:0] ? myVec_17 : _GEN_3770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3772 = 7'h12 == _myNewVec_99_T_3[6:0] ? myVec_18 : _GEN_3771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3773 = 7'h13 == _myNewVec_99_T_3[6:0] ? myVec_19 : _GEN_3772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3774 = 7'h14 == _myNewVec_99_T_3[6:0] ? myVec_20 : _GEN_3773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3775 = 7'h15 == _myNewVec_99_T_3[6:0] ? myVec_21 : _GEN_3774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3776 = 7'h16 == _myNewVec_99_T_3[6:0] ? myVec_22 : _GEN_3775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3777 = 7'h17 == _myNewVec_99_T_3[6:0] ? myVec_23 : _GEN_3776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3778 = 7'h18 == _myNewVec_99_T_3[6:0] ? myVec_24 : _GEN_3777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3779 = 7'h19 == _myNewVec_99_T_3[6:0] ? myVec_25 : _GEN_3778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3780 = 7'h1a == _myNewVec_99_T_3[6:0] ? myVec_26 : _GEN_3779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3781 = 7'h1b == _myNewVec_99_T_3[6:0] ? myVec_27 : _GEN_3780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3782 = 7'h1c == _myNewVec_99_T_3[6:0] ? myVec_28 : _GEN_3781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3783 = 7'h1d == _myNewVec_99_T_3[6:0] ? myVec_29 : _GEN_3782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3784 = 7'h1e == _myNewVec_99_T_3[6:0] ? myVec_30 : _GEN_3783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3785 = 7'h1f == _myNewVec_99_T_3[6:0] ? myVec_31 : _GEN_3784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3786 = 7'h20 == _myNewVec_99_T_3[6:0] ? myVec_32 : _GEN_3785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3787 = 7'h21 == _myNewVec_99_T_3[6:0] ? myVec_33 : _GEN_3786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3788 = 7'h22 == _myNewVec_99_T_3[6:0] ? myVec_34 : _GEN_3787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3789 = 7'h23 == _myNewVec_99_T_3[6:0] ? myVec_35 : _GEN_3788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3790 = 7'h24 == _myNewVec_99_T_3[6:0] ? myVec_36 : _GEN_3789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3791 = 7'h25 == _myNewVec_99_T_3[6:0] ? myVec_37 : _GEN_3790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3792 = 7'h26 == _myNewVec_99_T_3[6:0] ? myVec_38 : _GEN_3791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3793 = 7'h27 == _myNewVec_99_T_3[6:0] ? myVec_39 : _GEN_3792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3794 = 7'h28 == _myNewVec_99_T_3[6:0] ? myVec_40 : _GEN_3793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3795 = 7'h29 == _myNewVec_99_T_3[6:0] ? myVec_41 : _GEN_3794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3796 = 7'h2a == _myNewVec_99_T_3[6:0] ? myVec_42 : _GEN_3795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3797 = 7'h2b == _myNewVec_99_T_3[6:0] ? myVec_43 : _GEN_3796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3798 = 7'h2c == _myNewVec_99_T_3[6:0] ? myVec_44 : _GEN_3797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3799 = 7'h2d == _myNewVec_99_T_3[6:0] ? myVec_45 : _GEN_3798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3800 = 7'h2e == _myNewVec_99_T_3[6:0] ? myVec_46 : _GEN_3799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3801 = 7'h2f == _myNewVec_99_T_3[6:0] ? myVec_47 : _GEN_3800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3802 = 7'h30 == _myNewVec_99_T_3[6:0] ? myVec_48 : _GEN_3801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3803 = 7'h31 == _myNewVec_99_T_3[6:0] ? myVec_49 : _GEN_3802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3804 = 7'h32 == _myNewVec_99_T_3[6:0] ? myVec_50 : _GEN_3803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3805 = 7'h33 == _myNewVec_99_T_3[6:0] ? myVec_51 : _GEN_3804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3806 = 7'h34 == _myNewVec_99_T_3[6:0] ? myVec_52 : _GEN_3805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3807 = 7'h35 == _myNewVec_99_T_3[6:0] ? myVec_53 : _GEN_3806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3808 = 7'h36 == _myNewVec_99_T_3[6:0] ? myVec_54 : _GEN_3807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3809 = 7'h37 == _myNewVec_99_T_3[6:0] ? myVec_55 : _GEN_3808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3810 = 7'h38 == _myNewVec_99_T_3[6:0] ? myVec_56 : _GEN_3809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3811 = 7'h39 == _myNewVec_99_T_3[6:0] ? myVec_57 : _GEN_3810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3812 = 7'h3a == _myNewVec_99_T_3[6:0] ? myVec_58 : _GEN_3811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3813 = 7'h3b == _myNewVec_99_T_3[6:0] ? myVec_59 : _GEN_3812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3814 = 7'h3c == _myNewVec_99_T_3[6:0] ? myVec_60 : _GEN_3813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3815 = 7'h3d == _myNewVec_99_T_3[6:0] ? myVec_61 : _GEN_3814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3816 = 7'h3e == _myNewVec_99_T_3[6:0] ? myVec_62 : _GEN_3815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3817 = 7'h3f == _myNewVec_99_T_3[6:0] ? myVec_63 : _GEN_3816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3818 = 7'h40 == _myNewVec_99_T_3[6:0] ? myVec_64 : _GEN_3817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3819 = 7'h41 == _myNewVec_99_T_3[6:0] ? myVec_65 : _GEN_3818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3820 = 7'h42 == _myNewVec_99_T_3[6:0] ? myVec_66 : _GEN_3819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3821 = 7'h43 == _myNewVec_99_T_3[6:0] ? myVec_67 : _GEN_3820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3822 = 7'h44 == _myNewVec_99_T_3[6:0] ? myVec_68 : _GEN_3821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3823 = 7'h45 == _myNewVec_99_T_3[6:0] ? myVec_69 : _GEN_3822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3824 = 7'h46 == _myNewVec_99_T_3[6:0] ? myVec_70 : _GEN_3823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3825 = 7'h47 == _myNewVec_99_T_3[6:0] ? myVec_71 : _GEN_3824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3826 = 7'h48 == _myNewVec_99_T_3[6:0] ? myVec_72 : _GEN_3825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3827 = 7'h49 == _myNewVec_99_T_3[6:0] ? myVec_73 : _GEN_3826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3828 = 7'h4a == _myNewVec_99_T_3[6:0] ? myVec_74 : _GEN_3827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3829 = 7'h4b == _myNewVec_99_T_3[6:0] ? myVec_75 : _GEN_3828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3830 = 7'h4c == _myNewVec_99_T_3[6:0] ? myVec_76 : _GEN_3829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3831 = 7'h4d == _myNewVec_99_T_3[6:0] ? myVec_77 : _GEN_3830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3832 = 7'h4e == _myNewVec_99_T_3[6:0] ? myVec_78 : _GEN_3831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3833 = 7'h4f == _myNewVec_99_T_3[6:0] ? myVec_79 : _GEN_3832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3834 = 7'h50 == _myNewVec_99_T_3[6:0] ? myVec_80 : _GEN_3833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3835 = 7'h51 == _myNewVec_99_T_3[6:0] ? myVec_81 : _GEN_3834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3836 = 7'h52 == _myNewVec_99_T_3[6:0] ? myVec_82 : _GEN_3835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3837 = 7'h53 == _myNewVec_99_T_3[6:0] ? myVec_83 : _GEN_3836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3838 = 7'h54 == _myNewVec_99_T_3[6:0] ? myVec_84 : _GEN_3837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3839 = 7'h55 == _myNewVec_99_T_3[6:0] ? myVec_85 : _GEN_3838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3840 = 7'h56 == _myNewVec_99_T_3[6:0] ? myVec_86 : _GEN_3839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3841 = 7'h57 == _myNewVec_99_T_3[6:0] ? myVec_87 : _GEN_3840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3842 = 7'h58 == _myNewVec_99_T_3[6:0] ? myVec_88 : _GEN_3841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3843 = 7'h59 == _myNewVec_99_T_3[6:0] ? myVec_89 : _GEN_3842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3844 = 7'h5a == _myNewVec_99_T_3[6:0] ? myVec_90 : _GEN_3843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3845 = 7'h5b == _myNewVec_99_T_3[6:0] ? myVec_91 : _GEN_3844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3846 = 7'h5c == _myNewVec_99_T_3[6:0] ? myVec_92 : _GEN_3845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3847 = 7'h5d == _myNewVec_99_T_3[6:0] ? myVec_93 : _GEN_3846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3848 = 7'h5e == _myNewVec_99_T_3[6:0] ? myVec_94 : _GEN_3847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3849 = 7'h5f == _myNewVec_99_T_3[6:0] ? myVec_95 : _GEN_3848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3850 = 7'h60 == _myNewVec_99_T_3[6:0] ? myVec_96 : _GEN_3849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3851 = 7'h61 == _myNewVec_99_T_3[6:0] ? myVec_97 : _GEN_3850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3852 = 7'h62 == _myNewVec_99_T_3[6:0] ? myVec_98 : _GEN_3851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3853 = 7'h63 == _myNewVec_99_T_3[6:0] ? myVec_99 : _GEN_3852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3854 = 7'h64 == _myNewVec_99_T_3[6:0] ? myVec_100 : _GEN_3853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3855 = 7'h65 == _myNewVec_99_T_3[6:0] ? myVec_101 : _GEN_3854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3856 = 7'h66 == _myNewVec_99_T_3[6:0] ? myVec_102 : _GEN_3855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3857 = 7'h67 == _myNewVec_99_T_3[6:0] ? myVec_103 : _GEN_3856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3858 = 7'h68 == _myNewVec_99_T_3[6:0] ? myVec_104 : _GEN_3857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3859 = 7'h69 == _myNewVec_99_T_3[6:0] ? myVec_105 : _GEN_3858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3860 = 7'h6a == _myNewVec_99_T_3[6:0] ? myVec_106 : _GEN_3859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3861 = 7'h6b == _myNewVec_99_T_3[6:0] ? myVec_107 : _GEN_3860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3862 = 7'h6c == _myNewVec_99_T_3[6:0] ? myVec_108 : _GEN_3861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3863 = 7'h6d == _myNewVec_99_T_3[6:0] ? myVec_109 : _GEN_3862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3864 = 7'h6e == _myNewVec_99_T_3[6:0] ? myVec_110 : _GEN_3863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3865 = 7'h6f == _myNewVec_99_T_3[6:0] ? myVec_111 : _GEN_3864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3866 = 7'h70 == _myNewVec_99_T_3[6:0] ? myVec_112 : _GEN_3865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3867 = 7'h71 == _myNewVec_99_T_3[6:0] ? myVec_113 : _GEN_3866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3868 = 7'h72 == _myNewVec_99_T_3[6:0] ? myVec_114 : _GEN_3867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3869 = 7'h73 == _myNewVec_99_T_3[6:0] ? myVec_115 : _GEN_3868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3870 = 7'h74 == _myNewVec_99_T_3[6:0] ? myVec_116 : _GEN_3869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3871 = 7'h75 == _myNewVec_99_T_3[6:0] ? myVec_117 : _GEN_3870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3872 = 7'h76 == _myNewVec_99_T_3[6:0] ? myVec_118 : _GEN_3871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3873 = 7'h77 == _myNewVec_99_T_3[6:0] ? myVec_119 : _GEN_3872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3874 = 7'h78 == _myNewVec_99_T_3[6:0] ? myVec_120 : _GEN_3873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3875 = 7'h79 == _myNewVec_99_T_3[6:0] ? myVec_121 : _GEN_3874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3876 = 7'h7a == _myNewVec_99_T_3[6:0] ? myVec_122 : _GEN_3875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3877 = 7'h7b == _myNewVec_99_T_3[6:0] ? myVec_123 : _GEN_3876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3878 = 7'h7c == _myNewVec_99_T_3[6:0] ? myVec_124 : _GEN_3877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3879 = 7'h7d == _myNewVec_99_T_3[6:0] ? myVec_125 : _GEN_3878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3880 = 7'h7e == _myNewVec_99_T_3[6:0] ? myVec_126 : _GEN_3879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_99 = 7'h7f == _myNewVec_99_T_3[6:0] ? myVec_127 : _GEN_3880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_98_T_3 = _myNewVec_127_T_1 + 16'h1d; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3883 = 7'h1 == _myNewVec_98_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3884 = 7'h2 == _myNewVec_98_T_3[6:0] ? myVec_2 : _GEN_3883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3885 = 7'h3 == _myNewVec_98_T_3[6:0] ? myVec_3 : _GEN_3884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3886 = 7'h4 == _myNewVec_98_T_3[6:0] ? myVec_4 : _GEN_3885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3887 = 7'h5 == _myNewVec_98_T_3[6:0] ? myVec_5 : _GEN_3886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3888 = 7'h6 == _myNewVec_98_T_3[6:0] ? myVec_6 : _GEN_3887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3889 = 7'h7 == _myNewVec_98_T_3[6:0] ? myVec_7 : _GEN_3888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3890 = 7'h8 == _myNewVec_98_T_3[6:0] ? myVec_8 : _GEN_3889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3891 = 7'h9 == _myNewVec_98_T_3[6:0] ? myVec_9 : _GEN_3890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3892 = 7'ha == _myNewVec_98_T_3[6:0] ? myVec_10 : _GEN_3891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3893 = 7'hb == _myNewVec_98_T_3[6:0] ? myVec_11 : _GEN_3892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3894 = 7'hc == _myNewVec_98_T_3[6:0] ? myVec_12 : _GEN_3893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3895 = 7'hd == _myNewVec_98_T_3[6:0] ? myVec_13 : _GEN_3894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3896 = 7'he == _myNewVec_98_T_3[6:0] ? myVec_14 : _GEN_3895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3897 = 7'hf == _myNewVec_98_T_3[6:0] ? myVec_15 : _GEN_3896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3898 = 7'h10 == _myNewVec_98_T_3[6:0] ? myVec_16 : _GEN_3897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3899 = 7'h11 == _myNewVec_98_T_3[6:0] ? myVec_17 : _GEN_3898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3900 = 7'h12 == _myNewVec_98_T_3[6:0] ? myVec_18 : _GEN_3899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3901 = 7'h13 == _myNewVec_98_T_3[6:0] ? myVec_19 : _GEN_3900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3902 = 7'h14 == _myNewVec_98_T_3[6:0] ? myVec_20 : _GEN_3901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3903 = 7'h15 == _myNewVec_98_T_3[6:0] ? myVec_21 : _GEN_3902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3904 = 7'h16 == _myNewVec_98_T_3[6:0] ? myVec_22 : _GEN_3903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3905 = 7'h17 == _myNewVec_98_T_3[6:0] ? myVec_23 : _GEN_3904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3906 = 7'h18 == _myNewVec_98_T_3[6:0] ? myVec_24 : _GEN_3905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3907 = 7'h19 == _myNewVec_98_T_3[6:0] ? myVec_25 : _GEN_3906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3908 = 7'h1a == _myNewVec_98_T_3[6:0] ? myVec_26 : _GEN_3907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3909 = 7'h1b == _myNewVec_98_T_3[6:0] ? myVec_27 : _GEN_3908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3910 = 7'h1c == _myNewVec_98_T_3[6:0] ? myVec_28 : _GEN_3909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3911 = 7'h1d == _myNewVec_98_T_3[6:0] ? myVec_29 : _GEN_3910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3912 = 7'h1e == _myNewVec_98_T_3[6:0] ? myVec_30 : _GEN_3911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3913 = 7'h1f == _myNewVec_98_T_3[6:0] ? myVec_31 : _GEN_3912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3914 = 7'h20 == _myNewVec_98_T_3[6:0] ? myVec_32 : _GEN_3913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3915 = 7'h21 == _myNewVec_98_T_3[6:0] ? myVec_33 : _GEN_3914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3916 = 7'h22 == _myNewVec_98_T_3[6:0] ? myVec_34 : _GEN_3915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3917 = 7'h23 == _myNewVec_98_T_3[6:0] ? myVec_35 : _GEN_3916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3918 = 7'h24 == _myNewVec_98_T_3[6:0] ? myVec_36 : _GEN_3917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3919 = 7'h25 == _myNewVec_98_T_3[6:0] ? myVec_37 : _GEN_3918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3920 = 7'h26 == _myNewVec_98_T_3[6:0] ? myVec_38 : _GEN_3919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3921 = 7'h27 == _myNewVec_98_T_3[6:0] ? myVec_39 : _GEN_3920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3922 = 7'h28 == _myNewVec_98_T_3[6:0] ? myVec_40 : _GEN_3921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3923 = 7'h29 == _myNewVec_98_T_3[6:0] ? myVec_41 : _GEN_3922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3924 = 7'h2a == _myNewVec_98_T_3[6:0] ? myVec_42 : _GEN_3923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3925 = 7'h2b == _myNewVec_98_T_3[6:0] ? myVec_43 : _GEN_3924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3926 = 7'h2c == _myNewVec_98_T_3[6:0] ? myVec_44 : _GEN_3925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3927 = 7'h2d == _myNewVec_98_T_3[6:0] ? myVec_45 : _GEN_3926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3928 = 7'h2e == _myNewVec_98_T_3[6:0] ? myVec_46 : _GEN_3927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3929 = 7'h2f == _myNewVec_98_T_3[6:0] ? myVec_47 : _GEN_3928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3930 = 7'h30 == _myNewVec_98_T_3[6:0] ? myVec_48 : _GEN_3929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3931 = 7'h31 == _myNewVec_98_T_3[6:0] ? myVec_49 : _GEN_3930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3932 = 7'h32 == _myNewVec_98_T_3[6:0] ? myVec_50 : _GEN_3931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3933 = 7'h33 == _myNewVec_98_T_3[6:0] ? myVec_51 : _GEN_3932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3934 = 7'h34 == _myNewVec_98_T_3[6:0] ? myVec_52 : _GEN_3933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3935 = 7'h35 == _myNewVec_98_T_3[6:0] ? myVec_53 : _GEN_3934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3936 = 7'h36 == _myNewVec_98_T_3[6:0] ? myVec_54 : _GEN_3935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3937 = 7'h37 == _myNewVec_98_T_3[6:0] ? myVec_55 : _GEN_3936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3938 = 7'h38 == _myNewVec_98_T_3[6:0] ? myVec_56 : _GEN_3937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3939 = 7'h39 == _myNewVec_98_T_3[6:0] ? myVec_57 : _GEN_3938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3940 = 7'h3a == _myNewVec_98_T_3[6:0] ? myVec_58 : _GEN_3939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3941 = 7'h3b == _myNewVec_98_T_3[6:0] ? myVec_59 : _GEN_3940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3942 = 7'h3c == _myNewVec_98_T_3[6:0] ? myVec_60 : _GEN_3941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3943 = 7'h3d == _myNewVec_98_T_3[6:0] ? myVec_61 : _GEN_3942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3944 = 7'h3e == _myNewVec_98_T_3[6:0] ? myVec_62 : _GEN_3943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3945 = 7'h3f == _myNewVec_98_T_3[6:0] ? myVec_63 : _GEN_3944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3946 = 7'h40 == _myNewVec_98_T_3[6:0] ? myVec_64 : _GEN_3945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3947 = 7'h41 == _myNewVec_98_T_3[6:0] ? myVec_65 : _GEN_3946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3948 = 7'h42 == _myNewVec_98_T_3[6:0] ? myVec_66 : _GEN_3947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3949 = 7'h43 == _myNewVec_98_T_3[6:0] ? myVec_67 : _GEN_3948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3950 = 7'h44 == _myNewVec_98_T_3[6:0] ? myVec_68 : _GEN_3949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3951 = 7'h45 == _myNewVec_98_T_3[6:0] ? myVec_69 : _GEN_3950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3952 = 7'h46 == _myNewVec_98_T_3[6:0] ? myVec_70 : _GEN_3951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3953 = 7'h47 == _myNewVec_98_T_3[6:0] ? myVec_71 : _GEN_3952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3954 = 7'h48 == _myNewVec_98_T_3[6:0] ? myVec_72 : _GEN_3953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3955 = 7'h49 == _myNewVec_98_T_3[6:0] ? myVec_73 : _GEN_3954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3956 = 7'h4a == _myNewVec_98_T_3[6:0] ? myVec_74 : _GEN_3955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3957 = 7'h4b == _myNewVec_98_T_3[6:0] ? myVec_75 : _GEN_3956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3958 = 7'h4c == _myNewVec_98_T_3[6:0] ? myVec_76 : _GEN_3957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3959 = 7'h4d == _myNewVec_98_T_3[6:0] ? myVec_77 : _GEN_3958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3960 = 7'h4e == _myNewVec_98_T_3[6:0] ? myVec_78 : _GEN_3959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3961 = 7'h4f == _myNewVec_98_T_3[6:0] ? myVec_79 : _GEN_3960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3962 = 7'h50 == _myNewVec_98_T_3[6:0] ? myVec_80 : _GEN_3961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3963 = 7'h51 == _myNewVec_98_T_3[6:0] ? myVec_81 : _GEN_3962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3964 = 7'h52 == _myNewVec_98_T_3[6:0] ? myVec_82 : _GEN_3963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3965 = 7'h53 == _myNewVec_98_T_3[6:0] ? myVec_83 : _GEN_3964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3966 = 7'h54 == _myNewVec_98_T_3[6:0] ? myVec_84 : _GEN_3965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3967 = 7'h55 == _myNewVec_98_T_3[6:0] ? myVec_85 : _GEN_3966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3968 = 7'h56 == _myNewVec_98_T_3[6:0] ? myVec_86 : _GEN_3967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3969 = 7'h57 == _myNewVec_98_T_3[6:0] ? myVec_87 : _GEN_3968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3970 = 7'h58 == _myNewVec_98_T_3[6:0] ? myVec_88 : _GEN_3969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3971 = 7'h59 == _myNewVec_98_T_3[6:0] ? myVec_89 : _GEN_3970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3972 = 7'h5a == _myNewVec_98_T_3[6:0] ? myVec_90 : _GEN_3971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3973 = 7'h5b == _myNewVec_98_T_3[6:0] ? myVec_91 : _GEN_3972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3974 = 7'h5c == _myNewVec_98_T_3[6:0] ? myVec_92 : _GEN_3973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3975 = 7'h5d == _myNewVec_98_T_3[6:0] ? myVec_93 : _GEN_3974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3976 = 7'h5e == _myNewVec_98_T_3[6:0] ? myVec_94 : _GEN_3975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3977 = 7'h5f == _myNewVec_98_T_3[6:0] ? myVec_95 : _GEN_3976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3978 = 7'h60 == _myNewVec_98_T_3[6:0] ? myVec_96 : _GEN_3977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3979 = 7'h61 == _myNewVec_98_T_3[6:0] ? myVec_97 : _GEN_3978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3980 = 7'h62 == _myNewVec_98_T_3[6:0] ? myVec_98 : _GEN_3979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3981 = 7'h63 == _myNewVec_98_T_3[6:0] ? myVec_99 : _GEN_3980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3982 = 7'h64 == _myNewVec_98_T_3[6:0] ? myVec_100 : _GEN_3981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3983 = 7'h65 == _myNewVec_98_T_3[6:0] ? myVec_101 : _GEN_3982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3984 = 7'h66 == _myNewVec_98_T_3[6:0] ? myVec_102 : _GEN_3983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3985 = 7'h67 == _myNewVec_98_T_3[6:0] ? myVec_103 : _GEN_3984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3986 = 7'h68 == _myNewVec_98_T_3[6:0] ? myVec_104 : _GEN_3985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3987 = 7'h69 == _myNewVec_98_T_3[6:0] ? myVec_105 : _GEN_3986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3988 = 7'h6a == _myNewVec_98_T_3[6:0] ? myVec_106 : _GEN_3987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3989 = 7'h6b == _myNewVec_98_T_3[6:0] ? myVec_107 : _GEN_3988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3990 = 7'h6c == _myNewVec_98_T_3[6:0] ? myVec_108 : _GEN_3989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3991 = 7'h6d == _myNewVec_98_T_3[6:0] ? myVec_109 : _GEN_3990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3992 = 7'h6e == _myNewVec_98_T_3[6:0] ? myVec_110 : _GEN_3991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3993 = 7'h6f == _myNewVec_98_T_3[6:0] ? myVec_111 : _GEN_3992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3994 = 7'h70 == _myNewVec_98_T_3[6:0] ? myVec_112 : _GEN_3993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3995 = 7'h71 == _myNewVec_98_T_3[6:0] ? myVec_113 : _GEN_3994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3996 = 7'h72 == _myNewVec_98_T_3[6:0] ? myVec_114 : _GEN_3995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3997 = 7'h73 == _myNewVec_98_T_3[6:0] ? myVec_115 : _GEN_3996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3998 = 7'h74 == _myNewVec_98_T_3[6:0] ? myVec_116 : _GEN_3997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3999 = 7'h75 == _myNewVec_98_T_3[6:0] ? myVec_117 : _GEN_3998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4000 = 7'h76 == _myNewVec_98_T_3[6:0] ? myVec_118 : _GEN_3999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4001 = 7'h77 == _myNewVec_98_T_3[6:0] ? myVec_119 : _GEN_4000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4002 = 7'h78 == _myNewVec_98_T_3[6:0] ? myVec_120 : _GEN_4001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4003 = 7'h79 == _myNewVec_98_T_3[6:0] ? myVec_121 : _GEN_4002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4004 = 7'h7a == _myNewVec_98_T_3[6:0] ? myVec_122 : _GEN_4003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4005 = 7'h7b == _myNewVec_98_T_3[6:0] ? myVec_123 : _GEN_4004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4006 = 7'h7c == _myNewVec_98_T_3[6:0] ? myVec_124 : _GEN_4005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4007 = 7'h7d == _myNewVec_98_T_3[6:0] ? myVec_125 : _GEN_4006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4008 = 7'h7e == _myNewVec_98_T_3[6:0] ? myVec_126 : _GEN_4007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_98 = 7'h7f == _myNewVec_98_T_3[6:0] ? myVec_127 : _GEN_4008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_97_T_3 = _myNewVec_127_T_1 + 16'h1e; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_4011 = 7'h1 == _myNewVec_97_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4012 = 7'h2 == _myNewVec_97_T_3[6:0] ? myVec_2 : _GEN_4011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4013 = 7'h3 == _myNewVec_97_T_3[6:0] ? myVec_3 : _GEN_4012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4014 = 7'h4 == _myNewVec_97_T_3[6:0] ? myVec_4 : _GEN_4013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4015 = 7'h5 == _myNewVec_97_T_3[6:0] ? myVec_5 : _GEN_4014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4016 = 7'h6 == _myNewVec_97_T_3[6:0] ? myVec_6 : _GEN_4015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4017 = 7'h7 == _myNewVec_97_T_3[6:0] ? myVec_7 : _GEN_4016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4018 = 7'h8 == _myNewVec_97_T_3[6:0] ? myVec_8 : _GEN_4017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4019 = 7'h9 == _myNewVec_97_T_3[6:0] ? myVec_9 : _GEN_4018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4020 = 7'ha == _myNewVec_97_T_3[6:0] ? myVec_10 : _GEN_4019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4021 = 7'hb == _myNewVec_97_T_3[6:0] ? myVec_11 : _GEN_4020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4022 = 7'hc == _myNewVec_97_T_3[6:0] ? myVec_12 : _GEN_4021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4023 = 7'hd == _myNewVec_97_T_3[6:0] ? myVec_13 : _GEN_4022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4024 = 7'he == _myNewVec_97_T_3[6:0] ? myVec_14 : _GEN_4023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4025 = 7'hf == _myNewVec_97_T_3[6:0] ? myVec_15 : _GEN_4024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4026 = 7'h10 == _myNewVec_97_T_3[6:0] ? myVec_16 : _GEN_4025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4027 = 7'h11 == _myNewVec_97_T_3[6:0] ? myVec_17 : _GEN_4026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4028 = 7'h12 == _myNewVec_97_T_3[6:0] ? myVec_18 : _GEN_4027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4029 = 7'h13 == _myNewVec_97_T_3[6:0] ? myVec_19 : _GEN_4028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4030 = 7'h14 == _myNewVec_97_T_3[6:0] ? myVec_20 : _GEN_4029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4031 = 7'h15 == _myNewVec_97_T_3[6:0] ? myVec_21 : _GEN_4030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4032 = 7'h16 == _myNewVec_97_T_3[6:0] ? myVec_22 : _GEN_4031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4033 = 7'h17 == _myNewVec_97_T_3[6:0] ? myVec_23 : _GEN_4032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4034 = 7'h18 == _myNewVec_97_T_3[6:0] ? myVec_24 : _GEN_4033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4035 = 7'h19 == _myNewVec_97_T_3[6:0] ? myVec_25 : _GEN_4034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4036 = 7'h1a == _myNewVec_97_T_3[6:0] ? myVec_26 : _GEN_4035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4037 = 7'h1b == _myNewVec_97_T_3[6:0] ? myVec_27 : _GEN_4036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4038 = 7'h1c == _myNewVec_97_T_3[6:0] ? myVec_28 : _GEN_4037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4039 = 7'h1d == _myNewVec_97_T_3[6:0] ? myVec_29 : _GEN_4038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4040 = 7'h1e == _myNewVec_97_T_3[6:0] ? myVec_30 : _GEN_4039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4041 = 7'h1f == _myNewVec_97_T_3[6:0] ? myVec_31 : _GEN_4040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4042 = 7'h20 == _myNewVec_97_T_3[6:0] ? myVec_32 : _GEN_4041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4043 = 7'h21 == _myNewVec_97_T_3[6:0] ? myVec_33 : _GEN_4042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4044 = 7'h22 == _myNewVec_97_T_3[6:0] ? myVec_34 : _GEN_4043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4045 = 7'h23 == _myNewVec_97_T_3[6:0] ? myVec_35 : _GEN_4044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4046 = 7'h24 == _myNewVec_97_T_3[6:0] ? myVec_36 : _GEN_4045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4047 = 7'h25 == _myNewVec_97_T_3[6:0] ? myVec_37 : _GEN_4046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4048 = 7'h26 == _myNewVec_97_T_3[6:0] ? myVec_38 : _GEN_4047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4049 = 7'h27 == _myNewVec_97_T_3[6:0] ? myVec_39 : _GEN_4048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4050 = 7'h28 == _myNewVec_97_T_3[6:0] ? myVec_40 : _GEN_4049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4051 = 7'h29 == _myNewVec_97_T_3[6:0] ? myVec_41 : _GEN_4050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4052 = 7'h2a == _myNewVec_97_T_3[6:0] ? myVec_42 : _GEN_4051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4053 = 7'h2b == _myNewVec_97_T_3[6:0] ? myVec_43 : _GEN_4052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4054 = 7'h2c == _myNewVec_97_T_3[6:0] ? myVec_44 : _GEN_4053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4055 = 7'h2d == _myNewVec_97_T_3[6:0] ? myVec_45 : _GEN_4054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4056 = 7'h2e == _myNewVec_97_T_3[6:0] ? myVec_46 : _GEN_4055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4057 = 7'h2f == _myNewVec_97_T_3[6:0] ? myVec_47 : _GEN_4056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4058 = 7'h30 == _myNewVec_97_T_3[6:0] ? myVec_48 : _GEN_4057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4059 = 7'h31 == _myNewVec_97_T_3[6:0] ? myVec_49 : _GEN_4058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4060 = 7'h32 == _myNewVec_97_T_3[6:0] ? myVec_50 : _GEN_4059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4061 = 7'h33 == _myNewVec_97_T_3[6:0] ? myVec_51 : _GEN_4060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4062 = 7'h34 == _myNewVec_97_T_3[6:0] ? myVec_52 : _GEN_4061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4063 = 7'h35 == _myNewVec_97_T_3[6:0] ? myVec_53 : _GEN_4062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4064 = 7'h36 == _myNewVec_97_T_3[6:0] ? myVec_54 : _GEN_4063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4065 = 7'h37 == _myNewVec_97_T_3[6:0] ? myVec_55 : _GEN_4064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4066 = 7'h38 == _myNewVec_97_T_3[6:0] ? myVec_56 : _GEN_4065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4067 = 7'h39 == _myNewVec_97_T_3[6:0] ? myVec_57 : _GEN_4066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4068 = 7'h3a == _myNewVec_97_T_3[6:0] ? myVec_58 : _GEN_4067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4069 = 7'h3b == _myNewVec_97_T_3[6:0] ? myVec_59 : _GEN_4068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4070 = 7'h3c == _myNewVec_97_T_3[6:0] ? myVec_60 : _GEN_4069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4071 = 7'h3d == _myNewVec_97_T_3[6:0] ? myVec_61 : _GEN_4070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4072 = 7'h3e == _myNewVec_97_T_3[6:0] ? myVec_62 : _GEN_4071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4073 = 7'h3f == _myNewVec_97_T_3[6:0] ? myVec_63 : _GEN_4072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4074 = 7'h40 == _myNewVec_97_T_3[6:0] ? myVec_64 : _GEN_4073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4075 = 7'h41 == _myNewVec_97_T_3[6:0] ? myVec_65 : _GEN_4074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4076 = 7'h42 == _myNewVec_97_T_3[6:0] ? myVec_66 : _GEN_4075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4077 = 7'h43 == _myNewVec_97_T_3[6:0] ? myVec_67 : _GEN_4076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4078 = 7'h44 == _myNewVec_97_T_3[6:0] ? myVec_68 : _GEN_4077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4079 = 7'h45 == _myNewVec_97_T_3[6:0] ? myVec_69 : _GEN_4078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4080 = 7'h46 == _myNewVec_97_T_3[6:0] ? myVec_70 : _GEN_4079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4081 = 7'h47 == _myNewVec_97_T_3[6:0] ? myVec_71 : _GEN_4080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4082 = 7'h48 == _myNewVec_97_T_3[6:0] ? myVec_72 : _GEN_4081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4083 = 7'h49 == _myNewVec_97_T_3[6:0] ? myVec_73 : _GEN_4082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4084 = 7'h4a == _myNewVec_97_T_3[6:0] ? myVec_74 : _GEN_4083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4085 = 7'h4b == _myNewVec_97_T_3[6:0] ? myVec_75 : _GEN_4084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4086 = 7'h4c == _myNewVec_97_T_3[6:0] ? myVec_76 : _GEN_4085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4087 = 7'h4d == _myNewVec_97_T_3[6:0] ? myVec_77 : _GEN_4086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4088 = 7'h4e == _myNewVec_97_T_3[6:0] ? myVec_78 : _GEN_4087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4089 = 7'h4f == _myNewVec_97_T_3[6:0] ? myVec_79 : _GEN_4088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4090 = 7'h50 == _myNewVec_97_T_3[6:0] ? myVec_80 : _GEN_4089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4091 = 7'h51 == _myNewVec_97_T_3[6:0] ? myVec_81 : _GEN_4090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4092 = 7'h52 == _myNewVec_97_T_3[6:0] ? myVec_82 : _GEN_4091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4093 = 7'h53 == _myNewVec_97_T_3[6:0] ? myVec_83 : _GEN_4092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4094 = 7'h54 == _myNewVec_97_T_3[6:0] ? myVec_84 : _GEN_4093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4095 = 7'h55 == _myNewVec_97_T_3[6:0] ? myVec_85 : _GEN_4094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4096 = 7'h56 == _myNewVec_97_T_3[6:0] ? myVec_86 : _GEN_4095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4097 = 7'h57 == _myNewVec_97_T_3[6:0] ? myVec_87 : _GEN_4096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4098 = 7'h58 == _myNewVec_97_T_3[6:0] ? myVec_88 : _GEN_4097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4099 = 7'h59 == _myNewVec_97_T_3[6:0] ? myVec_89 : _GEN_4098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4100 = 7'h5a == _myNewVec_97_T_3[6:0] ? myVec_90 : _GEN_4099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4101 = 7'h5b == _myNewVec_97_T_3[6:0] ? myVec_91 : _GEN_4100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4102 = 7'h5c == _myNewVec_97_T_3[6:0] ? myVec_92 : _GEN_4101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4103 = 7'h5d == _myNewVec_97_T_3[6:0] ? myVec_93 : _GEN_4102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4104 = 7'h5e == _myNewVec_97_T_3[6:0] ? myVec_94 : _GEN_4103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4105 = 7'h5f == _myNewVec_97_T_3[6:0] ? myVec_95 : _GEN_4104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4106 = 7'h60 == _myNewVec_97_T_3[6:0] ? myVec_96 : _GEN_4105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4107 = 7'h61 == _myNewVec_97_T_3[6:0] ? myVec_97 : _GEN_4106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4108 = 7'h62 == _myNewVec_97_T_3[6:0] ? myVec_98 : _GEN_4107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4109 = 7'h63 == _myNewVec_97_T_3[6:0] ? myVec_99 : _GEN_4108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4110 = 7'h64 == _myNewVec_97_T_3[6:0] ? myVec_100 : _GEN_4109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4111 = 7'h65 == _myNewVec_97_T_3[6:0] ? myVec_101 : _GEN_4110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4112 = 7'h66 == _myNewVec_97_T_3[6:0] ? myVec_102 : _GEN_4111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4113 = 7'h67 == _myNewVec_97_T_3[6:0] ? myVec_103 : _GEN_4112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4114 = 7'h68 == _myNewVec_97_T_3[6:0] ? myVec_104 : _GEN_4113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4115 = 7'h69 == _myNewVec_97_T_3[6:0] ? myVec_105 : _GEN_4114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4116 = 7'h6a == _myNewVec_97_T_3[6:0] ? myVec_106 : _GEN_4115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4117 = 7'h6b == _myNewVec_97_T_3[6:0] ? myVec_107 : _GEN_4116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4118 = 7'h6c == _myNewVec_97_T_3[6:0] ? myVec_108 : _GEN_4117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4119 = 7'h6d == _myNewVec_97_T_3[6:0] ? myVec_109 : _GEN_4118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4120 = 7'h6e == _myNewVec_97_T_3[6:0] ? myVec_110 : _GEN_4119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4121 = 7'h6f == _myNewVec_97_T_3[6:0] ? myVec_111 : _GEN_4120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4122 = 7'h70 == _myNewVec_97_T_3[6:0] ? myVec_112 : _GEN_4121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4123 = 7'h71 == _myNewVec_97_T_3[6:0] ? myVec_113 : _GEN_4122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4124 = 7'h72 == _myNewVec_97_T_3[6:0] ? myVec_114 : _GEN_4123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4125 = 7'h73 == _myNewVec_97_T_3[6:0] ? myVec_115 : _GEN_4124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4126 = 7'h74 == _myNewVec_97_T_3[6:0] ? myVec_116 : _GEN_4125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4127 = 7'h75 == _myNewVec_97_T_3[6:0] ? myVec_117 : _GEN_4126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4128 = 7'h76 == _myNewVec_97_T_3[6:0] ? myVec_118 : _GEN_4127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4129 = 7'h77 == _myNewVec_97_T_3[6:0] ? myVec_119 : _GEN_4128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4130 = 7'h78 == _myNewVec_97_T_3[6:0] ? myVec_120 : _GEN_4129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4131 = 7'h79 == _myNewVec_97_T_3[6:0] ? myVec_121 : _GEN_4130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4132 = 7'h7a == _myNewVec_97_T_3[6:0] ? myVec_122 : _GEN_4131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4133 = 7'h7b == _myNewVec_97_T_3[6:0] ? myVec_123 : _GEN_4132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4134 = 7'h7c == _myNewVec_97_T_3[6:0] ? myVec_124 : _GEN_4133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4135 = 7'h7d == _myNewVec_97_T_3[6:0] ? myVec_125 : _GEN_4134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4136 = 7'h7e == _myNewVec_97_T_3[6:0] ? myVec_126 : _GEN_4135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_97 = 7'h7f == _myNewVec_97_T_3[6:0] ? myVec_127 : _GEN_4136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_96_T_3 = _myNewVec_127_T_1 + 16'h1f; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_4139 = 7'h1 == _myNewVec_96_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4140 = 7'h2 == _myNewVec_96_T_3[6:0] ? myVec_2 : _GEN_4139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4141 = 7'h3 == _myNewVec_96_T_3[6:0] ? myVec_3 : _GEN_4140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4142 = 7'h4 == _myNewVec_96_T_3[6:0] ? myVec_4 : _GEN_4141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4143 = 7'h5 == _myNewVec_96_T_3[6:0] ? myVec_5 : _GEN_4142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4144 = 7'h6 == _myNewVec_96_T_3[6:0] ? myVec_6 : _GEN_4143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4145 = 7'h7 == _myNewVec_96_T_3[6:0] ? myVec_7 : _GEN_4144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4146 = 7'h8 == _myNewVec_96_T_3[6:0] ? myVec_8 : _GEN_4145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4147 = 7'h9 == _myNewVec_96_T_3[6:0] ? myVec_9 : _GEN_4146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4148 = 7'ha == _myNewVec_96_T_3[6:0] ? myVec_10 : _GEN_4147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4149 = 7'hb == _myNewVec_96_T_3[6:0] ? myVec_11 : _GEN_4148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4150 = 7'hc == _myNewVec_96_T_3[6:0] ? myVec_12 : _GEN_4149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4151 = 7'hd == _myNewVec_96_T_3[6:0] ? myVec_13 : _GEN_4150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4152 = 7'he == _myNewVec_96_T_3[6:0] ? myVec_14 : _GEN_4151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4153 = 7'hf == _myNewVec_96_T_3[6:0] ? myVec_15 : _GEN_4152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4154 = 7'h10 == _myNewVec_96_T_3[6:0] ? myVec_16 : _GEN_4153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4155 = 7'h11 == _myNewVec_96_T_3[6:0] ? myVec_17 : _GEN_4154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4156 = 7'h12 == _myNewVec_96_T_3[6:0] ? myVec_18 : _GEN_4155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4157 = 7'h13 == _myNewVec_96_T_3[6:0] ? myVec_19 : _GEN_4156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4158 = 7'h14 == _myNewVec_96_T_3[6:0] ? myVec_20 : _GEN_4157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4159 = 7'h15 == _myNewVec_96_T_3[6:0] ? myVec_21 : _GEN_4158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4160 = 7'h16 == _myNewVec_96_T_3[6:0] ? myVec_22 : _GEN_4159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4161 = 7'h17 == _myNewVec_96_T_3[6:0] ? myVec_23 : _GEN_4160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4162 = 7'h18 == _myNewVec_96_T_3[6:0] ? myVec_24 : _GEN_4161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4163 = 7'h19 == _myNewVec_96_T_3[6:0] ? myVec_25 : _GEN_4162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4164 = 7'h1a == _myNewVec_96_T_3[6:0] ? myVec_26 : _GEN_4163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4165 = 7'h1b == _myNewVec_96_T_3[6:0] ? myVec_27 : _GEN_4164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4166 = 7'h1c == _myNewVec_96_T_3[6:0] ? myVec_28 : _GEN_4165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4167 = 7'h1d == _myNewVec_96_T_3[6:0] ? myVec_29 : _GEN_4166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4168 = 7'h1e == _myNewVec_96_T_3[6:0] ? myVec_30 : _GEN_4167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4169 = 7'h1f == _myNewVec_96_T_3[6:0] ? myVec_31 : _GEN_4168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4170 = 7'h20 == _myNewVec_96_T_3[6:0] ? myVec_32 : _GEN_4169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4171 = 7'h21 == _myNewVec_96_T_3[6:0] ? myVec_33 : _GEN_4170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4172 = 7'h22 == _myNewVec_96_T_3[6:0] ? myVec_34 : _GEN_4171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4173 = 7'h23 == _myNewVec_96_T_3[6:0] ? myVec_35 : _GEN_4172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4174 = 7'h24 == _myNewVec_96_T_3[6:0] ? myVec_36 : _GEN_4173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4175 = 7'h25 == _myNewVec_96_T_3[6:0] ? myVec_37 : _GEN_4174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4176 = 7'h26 == _myNewVec_96_T_3[6:0] ? myVec_38 : _GEN_4175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4177 = 7'h27 == _myNewVec_96_T_3[6:0] ? myVec_39 : _GEN_4176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4178 = 7'h28 == _myNewVec_96_T_3[6:0] ? myVec_40 : _GEN_4177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4179 = 7'h29 == _myNewVec_96_T_3[6:0] ? myVec_41 : _GEN_4178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4180 = 7'h2a == _myNewVec_96_T_3[6:0] ? myVec_42 : _GEN_4179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4181 = 7'h2b == _myNewVec_96_T_3[6:0] ? myVec_43 : _GEN_4180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4182 = 7'h2c == _myNewVec_96_T_3[6:0] ? myVec_44 : _GEN_4181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4183 = 7'h2d == _myNewVec_96_T_3[6:0] ? myVec_45 : _GEN_4182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4184 = 7'h2e == _myNewVec_96_T_3[6:0] ? myVec_46 : _GEN_4183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4185 = 7'h2f == _myNewVec_96_T_3[6:0] ? myVec_47 : _GEN_4184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4186 = 7'h30 == _myNewVec_96_T_3[6:0] ? myVec_48 : _GEN_4185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4187 = 7'h31 == _myNewVec_96_T_3[6:0] ? myVec_49 : _GEN_4186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4188 = 7'h32 == _myNewVec_96_T_3[6:0] ? myVec_50 : _GEN_4187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4189 = 7'h33 == _myNewVec_96_T_3[6:0] ? myVec_51 : _GEN_4188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4190 = 7'h34 == _myNewVec_96_T_3[6:0] ? myVec_52 : _GEN_4189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4191 = 7'h35 == _myNewVec_96_T_3[6:0] ? myVec_53 : _GEN_4190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4192 = 7'h36 == _myNewVec_96_T_3[6:0] ? myVec_54 : _GEN_4191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4193 = 7'h37 == _myNewVec_96_T_3[6:0] ? myVec_55 : _GEN_4192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4194 = 7'h38 == _myNewVec_96_T_3[6:0] ? myVec_56 : _GEN_4193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4195 = 7'h39 == _myNewVec_96_T_3[6:0] ? myVec_57 : _GEN_4194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4196 = 7'h3a == _myNewVec_96_T_3[6:0] ? myVec_58 : _GEN_4195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4197 = 7'h3b == _myNewVec_96_T_3[6:0] ? myVec_59 : _GEN_4196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4198 = 7'h3c == _myNewVec_96_T_3[6:0] ? myVec_60 : _GEN_4197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4199 = 7'h3d == _myNewVec_96_T_3[6:0] ? myVec_61 : _GEN_4198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4200 = 7'h3e == _myNewVec_96_T_3[6:0] ? myVec_62 : _GEN_4199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4201 = 7'h3f == _myNewVec_96_T_3[6:0] ? myVec_63 : _GEN_4200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4202 = 7'h40 == _myNewVec_96_T_3[6:0] ? myVec_64 : _GEN_4201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4203 = 7'h41 == _myNewVec_96_T_3[6:0] ? myVec_65 : _GEN_4202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4204 = 7'h42 == _myNewVec_96_T_3[6:0] ? myVec_66 : _GEN_4203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4205 = 7'h43 == _myNewVec_96_T_3[6:0] ? myVec_67 : _GEN_4204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4206 = 7'h44 == _myNewVec_96_T_3[6:0] ? myVec_68 : _GEN_4205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4207 = 7'h45 == _myNewVec_96_T_3[6:0] ? myVec_69 : _GEN_4206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4208 = 7'h46 == _myNewVec_96_T_3[6:0] ? myVec_70 : _GEN_4207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4209 = 7'h47 == _myNewVec_96_T_3[6:0] ? myVec_71 : _GEN_4208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4210 = 7'h48 == _myNewVec_96_T_3[6:0] ? myVec_72 : _GEN_4209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4211 = 7'h49 == _myNewVec_96_T_3[6:0] ? myVec_73 : _GEN_4210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4212 = 7'h4a == _myNewVec_96_T_3[6:0] ? myVec_74 : _GEN_4211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4213 = 7'h4b == _myNewVec_96_T_3[6:0] ? myVec_75 : _GEN_4212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4214 = 7'h4c == _myNewVec_96_T_3[6:0] ? myVec_76 : _GEN_4213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4215 = 7'h4d == _myNewVec_96_T_3[6:0] ? myVec_77 : _GEN_4214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4216 = 7'h4e == _myNewVec_96_T_3[6:0] ? myVec_78 : _GEN_4215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4217 = 7'h4f == _myNewVec_96_T_3[6:0] ? myVec_79 : _GEN_4216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4218 = 7'h50 == _myNewVec_96_T_3[6:0] ? myVec_80 : _GEN_4217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4219 = 7'h51 == _myNewVec_96_T_3[6:0] ? myVec_81 : _GEN_4218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4220 = 7'h52 == _myNewVec_96_T_3[6:0] ? myVec_82 : _GEN_4219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4221 = 7'h53 == _myNewVec_96_T_3[6:0] ? myVec_83 : _GEN_4220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4222 = 7'h54 == _myNewVec_96_T_3[6:0] ? myVec_84 : _GEN_4221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4223 = 7'h55 == _myNewVec_96_T_3[6:0] ? myVec_85 : _GEN_4222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4224 = 7'h56 == _myNewVec_96_T_3[6:0] ? myVec_86 : _GEN_4223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4225 = 7'h57 == _myNewVec_96_T_3[6:0] ? myVec_87 : _GEN_4224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4226 = 7'h58 == _myNewVec_96_T_3[6:0] ? myVec_88 : _GEN_4225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4227 = 7'h59 == _myNewVec_96_T_3[6:0] ? myVec_89 : _GEN_4226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4228 = 7'h5a == _myNewVec_96_T_3[6:0] ? myVec_90 : _GEN_4227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4229 = 7'h5b == _myNewVec_96_T_3[6:0] ? myVec_91 : _GEN_4228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4230 = 7'h5c == _myNewVec_96_T_3[6:0] ? myVec_92 : _GEN_4229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4231 = 7'h5d == _myNewVec_96_T_3[6:0] ? myVec_93 : _GEN_4230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4232 = 7'h5e == _myNewVec_96_T_3[6:0] ? myVec_94 : _GEN_4231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4233 = 7'h5f == _myNewVec_96_T_3[6:0] ? myVec_95 : _GEN_4232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4234 = 7'h60 == _myNewVec_96_T_3[6:0] ? myVec_96 : _GEN_4233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4235 = 7'h61 == _myNewVec_96_T_3[6:0] ? myVec_97 : _GEN_4234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4236 = 7'h62 == _myNewVec_96_T_3[6:0] ? myVec_98 : _GEN_4235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4237 = 7'h63 == _myNewVec_96_T_3[6:0] ? myVec_99 : _GEN_4236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4238 = 7'h64 == _myNewVec_96_T_3[6:0] ? myVec_100 : _GEN_4237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4239 = 7'h65 == _myNewVec_96_T_3[6:0] ? myVec_101 : _GEN_4238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4240 = 7'h66 == _myNewVec_96_T_3[6:0] ? myVec_102 : _GEN_4239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4241 = 7'h67 == _myNewVec_96_T_3[6:0] ? myVec_103 : _GEN_4240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4242 = 7'h68 == _myNewVec_96_T_3[6:0] ? myVec_104 : _GEN_4241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4243 = 7'h69 == _myNewVec_96_T_3[6:0] ? myVec_105 : _GEN_4242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4244 = 7'h6a == _myNewVec_96_T_3[6:0] ? myVec_106 : _GEN_4243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4245 = 7'h6b == _myNewVec_96_T_3[6:0] ? myVec_107 : _GEN_4244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4246 = 7'h6c == _myNewVec_96_T_3[6:0] ? myVec_108 : _GEN_4245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4247 = 7'h6d == _myNewVec_96_T_3[6:0] ? myVec_109 : _GEN_4246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4248 = 7'h6e == _myNewVec_96_T_3[6:0] ? myVec_110 : _GEN_4247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4249 = 7'h6f == _myNewVec_96_T_3[6:0] ? myVec_111 : _GEN_4248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4250 = 7'h70 == _myNewVec_96_T_3[6:0] ? myVec_112 : _GEN_4249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4251 = 7'h71 == _myNewVec_96_T_3[6:0] ? myVec_113 : _GEN_4250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4252 = 7'h72 == _myNewVec_96_T_3[6:0] ? myVec_114 : _GEN_4251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4253 = 7'h73 == _myNewVec_96_T_3[6:0] ? myVec_115 : _GEN_4252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4254 = 7'h74 == _myNewVec_96_T_3[6:0] ? myVec_116 : _GEN_4253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4255 = 7'h75 == _myNewVec_96_T_3[6:0] ? myVec_117 : _GEN_4254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4256 = 7'h76 == _myNewVec_96_T_3[6:0] ? myVec_118 : _GEN_4255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4257 = 7'h77 == _myNewVec_96_T_3[6:0] ? myVec_119 : _GEN_4256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4258 = 7'h78 == _myNewVec_96_T_3[6:0] ? myVec_120 : _GEN_4257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4259 = 7'h79 == _myNewVec_96_T_3[6:0] ? myVec_121 : _GEN_4258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4260 = 7'h7a == _myNewVec_96_T_3[6:0] ? myVec_122 : _GEN_4259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4261 = 7'h7b == _myNewVec_96_T_3[6:0] ? myVec_123 : _GEN_4260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4262 = 7'h7c == _myNewVec_96_T_3[6:0] ? myVec_124 : _GEN_4261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4263 = 7'h7d == _myNewVec_96_T_3[6:0] ? myVec_125 : _GEN_4262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4264 = 7'h7e == _myNewVec_96_T_3[6:0] ? myVec_126 : _GEN_4263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_96 = 7'h7f == _myNewVec_96_T_3[6:0] ? myVec_127 : _GEN_4264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [255:0] myNewWire_hi_hi_lo_lo = {myNewVec_103,myNewVec_102,myNewVec_101,myNewVec_100,myNewVec_99,myNewVec_98,
    myNewVec_97,myNewVec_96}; // @[hh_datapath_chisel.scala 238:27]
  wire [511:0] myNewWire_hi_hi_lo = {myNewVec_111,myNewVec_110,myNewVec_109,myNewVec_108,myNewVec_107,myNewVec_106,
    myNewVec_105,myNewVec_104,myNewWire_hi_hi_lo_lo}; // @[hh_datapath_chisel.scala 238:27]
  wire [1023:0] myNewWire_hi_hi = {myNewVec_127,myNewVec_126,myNewVec_125,myNewVec_124,myNewVec_123,myNewVec_122,
    myNewVec_121,myNewVec_120,myNewWire_hi_hi_hi_lo,myNewWire_hi_hi_lo}; // @[hh_datapath_chisel.scala 238:27]
  wire [15:0] _myNewVec_95_T_3 = _myNewVec_127_T_1 + 16'h20; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_4267 = 7'h1 == _myNewVec_95_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4268 = 7'h2 == _myNewVec_95_T_3[6:0] ? myVec_2 : _GEN_4267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4269 = 7'h3 == _myNewVec_95_T_3[6:0] ? myVec_3 : _GEN_4268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4270 = 7'h4 == _myNewVec_95_T_3[6:0] ? myVec_4 : _GEN_4269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4271 = 7'h5 == _myNewVec_95_T_3[6:0] ? myVec_5 : _GEN_4270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4272 = 7'h6 == _myNewVec_95_T_3[6:0] ? myVec_6 : _GEN_4271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4273 = 7'h7 == _myNewVec_95_T_3[6:0] ? myVec_7 : _GEN_4272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4274 = 7'h8 == _myNewVec_95_T_3[6:0] ? myVec_8 : _GEN_4273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4275 = 7'h9 == _myNewVec_95_T_3[6:0] ? myVec_9 : _GEN_4274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4276 = 7'ha == _myNewVec_95_T_3[6:0] ? myVec_10 : _GEN_4275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4277 = 7'hb == _myNewVec_95_T_3[6:0] ? myVec_11 : _GEN_4276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4278 = 7'hc == _myNewVec_95_T_3[6:0] ? myVec_12 : _GEN_4277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4279 = 7'hd == _myNewVec_95_T_3[6:0] ? myVec_13 : _GEN_4278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4280 = 7'he == _myNewVec_95_T_3[6:0] ? myVec_14 : _GEN_4279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4281 = 7'hf == _myNewVec_95_T_3[6:0] ? myVec_15 : _GEN_4280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4282 = 7'h10 == _myNewVec_95_T_3[6:0] ? myVec_16 : _GEN_4281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4283 = 7'h11 == _myNewVec_95_T_3[6:0] ? myVec_17 : _GEN_4282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4284 = 7'h12 == _myNewVec_95_T_3[6:0] ? myVec_18 : _GEN_4283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4285 = 7'h13 == _myNewVec_95_T_3[6:0] ? myVec_19 : _GEN_4284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4286 = 7'h14 == _myNewVec_95_T_3[6:0] ? myVec_20 : _GEN_4285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4287 = 7'h15 == _myNewVec_95_T_3[6:0] ? myVec_21 : _GEN_4286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4288 = 7'h16 == _myNewVec_95_T_3[6:0] ? myVec_22 : _GEN_4287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4289 = 7'h17 == _myNewVec_95_T_3[6:0] ? myVec_23 : _GEN_4288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4290 = 7'h18 == _myNewVec_95_T_3[6:0] ? myVec_24 : _GEN_4289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4291 = 7'h19 == _myNewVec_95_T_3[6:0] ? myVec_25 : _GEN_4290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4292 = 7'h1a == _myNewVec_95_T_3[6:0] ? myVec_26 : _GEN_4291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4293 = 7'h1b == _myNewVec_95_T_3[6:0] ? myVec_27 : _GEN_4292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4294 = 7'h1c == _myNewVec_95_T_3[6:0] ? myVec_28 : _GEN_4293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4295 = 7'h1d == _myNewVec_95_T_3[6:0] ? myVec_29 : _GEN_4294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4296 = 7'h1e == _myNewVec_95_T_3[6:0] ? myVec_30 : _GEN_4295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4297 = 7'h1f == _myNewVec_95_T_3[6:0] ? myVec_31 : _GEN_4296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4298 = 7'h20 == _myNewVec_95_T_3[6:0] ? myVec_32 : _GEN_4297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4299 = 7'h21 == _myNewVec_95_T_3[6:0] ? myVec_33 : _GEN_4298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4300 = 7'h22 == _myNewVec_95_T_3[6:0] ? myVec_34 : _GEN_4299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4301 = 7'h23 == _myNewVec_95_T_3[6:0] ? myVec_35 : _GEN_4300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4302 = 7'h24 == _myNewVec_95_T_3[6:0] ? myVec_36 : _GEN_4301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4303 = 7'h25 == _myNewVec_95_T_3[6:0] ? myVec_37 : _GEN_4302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4304 = 7'h26 == _myNewVec_95_T_3[6:0] ? myVec_38 : _GEN_4303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4305 = 7'h27 == _myNewVec_95_T_3[6:0] ? myVec_39 : _GEN_4304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4306 = 7'h28 == _myNewVec_95_T_3[6:0] ? myVec_40 : _GEN_4305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4307 = 7'h29 == _myNewVec_95_T_3[6:0] ? myVec_41 : _GEN_4306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4308 = 7'h2a == _myNewVec_95_T_3[6:0] ? myVec_42 : _GEN_4307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4309 = 7'h2b == _myNewVec_95_T_3[6:0] ? myVec_43 : _GEN_4308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4310 = 7'h2c == _myNewVec_95_T_3[6:0] ? myVec_44 : _GEN_4309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4311 = 7'h2d == _myNewVec_95_T_3[6:0] ? myVec_45 : _GEN_4310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4312 = 7'h2e == _myNewVec_95_T_3[6:0] ? myVec_46 : _GEN_4311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4313 = 7'h2f == _myNewVec_95_T_3[6:0] ? myVec_47 : _GEN_4312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4314 = 7'h30 == _myNewVec_95_T_3[6:0] ? myVec_48 : _GEN_4313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4315 = 7'h31 == _myNewVec_95_T_3[6:0] ? myVec_49 : _GEN_4314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4316 = 7'h32 == _myNewVec_95_T_3[6:0] ? myVec_50 : _GEN_4315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4317 = 7'h33 == _myNewVec_95_T_3[6:0] ? myVec_51 : _GEN_4316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4318 = 7'h34 == _myNewVec_95_T_3[6:0] ? myVec_52 : _GEN_4317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4319 = 7'h35 == _myNewVec_95_T_3[6:0] ? myVec_53 : _GEN_4318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4320 = 7'h36 == _myNewVec_95_T_3[6:0] ? myVec_54 : _GEN_4319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4321 = 7'h37 == _myNewVec_95_T_3[6:0] ? myVec_55 : _GEN_4320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4322 = 7'h38 == _myNewVec_95_T_3[6:0] ? myVec_56 : _GEN_4321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4323 = 7'h39 == _myNewVec_95_T_3[6:0] ? myVec_57 : _GEN_4322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4324 = 7'h3a == _myNewVec_95_T_3[6:0] ? myVec_58 : _GEN_4323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4325 = 7'h3b == _myNewVec_95_T_3[6:0] ? myVec_59 : _GEN_4324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4326 = 7'h3c == _myNewVec_95_T_3[6:0] ? myVec_60 : _GEN_4325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4327 = 7'h3d == _myNewVec_95_T_3[6:0] ? myVec_61 : _GEN_4326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4328 = 7'h3e == _myNewVec_95_T_3[6:0] ? myVec_62 : _GEN_4327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4329 = 7'h3f == _myNewVec_95_T_3[6:0] ? myVec_63 : _GEN_4328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4330 = 7'h40 == _myNewVec_95_T_3[6:0] ? myVec_64 : _GEN_4329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4331 = 7'h41 == _myNewVec_95_T_3[6:0] ? myVec_65 : _GEN_4330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4332 = 7'h42 == _myNewVec_95_T_3[6:0] ? myVec_66 : _GEN_4331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4333 = 7'h43 == _myNewVec_95_T_3[6:0] ? myVec_67 : _GEN_4332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4334 = 7'h44 == _myNewVec_95_T_3[6:0] ? myVec_68 : _GEN_4333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4335 = 7'h45 == _myNewVec_95_T_3[6:0] ? myVec_69 : _GEN_4334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4336 = 7'h46 == _myNewVec_95_T_3[6:0] ? myVec_70 : _GEN_4335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4337 = 7'h47 == _myNewVec_95_T_3[6:0] ? myVec_71 : _GEN_4336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4338 = 7'h48 == _myNewVec_95_T_3[6:0] ? myVec_72 : _GEN_4337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4339 = 7'h49 == _myNewVec_95_T_3[6:0] ? myVec_73 : _GEN_4338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4340 = 7'h4a == _myNewVec_95_T_3[6:0] ? myVec_74 : _GEN_4339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4341 = 7'h4b == _myNewVec_95_T_3[6:0] ? myVec_75 : _GEN_4340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4342 = 7'h4c == _myNewVec_95_T_3[6:0] ? myVec_76 : _GEN_4341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4343 = 7'h4d == _myNewVec_95_T_3[6:0] ? myVec_77 : _GEN_4342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4344 = 7'h4e == _myNewVec_95_T_3[6:0] ? myVec_78 : _GEN_4343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4345 = 7'h4f == _myNewVec_95_T_3[6:0] ? myVec_79 : _GEN_4344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4346 = 7'h50 == _myNewVec_95_T_3[6:0] ? myVec_80 : _GEN_4345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4347 = 7'h51 == _myNewVec_95_T_3[6:0] ? myVec_81 : _GEN_4346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4348 = 7'h52 == _myNewVec_95_T_3[6:0] ? myVec_82 : _GEN_4347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4349 = 7'h53 == _myNewVec_95_T_3[6:0] ? myVec_83 : _GEN_4348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4350 = 7'h54 == _myNewVec_95_T_3[6:0] ? myVec_84 : _GEN_4349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4351 = 7'h55 == _myNewVec_95_T_3[6:0] ? myVec_85 : _GEN_4350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4352 = 7'h56 == _myNewVec_95_T_3[6:0] ? myVec_86 : _GEN_4351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4353 = 7'h57 == _myNewVec_95_T_3[6:0] ? myVec_87 : _GEN_4352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4354 = 7'h58 == _myNewVec_95_T_3[6:0] ? myVec_88 : _GEN_4353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4355 = 7'h59 == _myNewVec_95_T_3[6:0] ? myVec_89 : _GEN_4354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4356 = 7'h5a == _myNewVec_95_T_3[6:0] ? myVec_90 : _GEN_4355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4357 = 7'h5b == _myNewVec_95_T_3[6:0] ? myVec_91 : _GEN_4356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4358 = 7'h5c == _myNewVec_95_T_3[6:0] ? myVec_92 : _GEN_4357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4359 = 7'h5d == _myNewVec_95_T_3[6:0] ? myVec_93 : _GEN_4358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4360 = 7'h5e == _myNewVec_95_T_3[6:0] ? myVec_94 : _GEN_4359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4361 = 7'h5f == _myNewVec_95_T_3[6:0] ? myVec_95 : _GEN_4360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4362 = 7'h60 == _myNewVec_95_T_3[6:0] ? myVec_96 : _GEN_4361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4363 = 7'h61 == _myNewVec_95_T_3[6:0] ? myVec_97 : _GEN_4362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4364 = 7'h62 == _myNewVec_95_T_3[6:0] ? myVec_98 : _GEN_4363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4365 = 7'h63 == _myNewVec_95_T_3[6:0] ? myVec_99 : _GEN_4364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4366 = 7'h64 == _myNewVec_95_T_3[6:0] ? myVec_100 : _GEN_4365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4367 = 7'h65 == _myNewVec_95_T_3[6:0] ? myVec_101 : _GEN_4366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4368 = 7'h66 == _myNewVec_95_T_3[6:0] ? myVec_102 : _GEN_4367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4369 = 7'h67 == _myNewVec_95_T_3[6:0] ? myVec_103 : _GEN_4368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4370 = 7'h68 == _myNewVec_95_T_3[6:0] ? myVec_104 : _GEN_4369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4371 = 7'h69 == _myNewVec_95_T_3[6:0] ? myVec_105 : _GEN_4370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4372 = 7'h6a == _myNewVec_95_T_3[6:0] ? myVec_106 : _GEN_4371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4373 = 7'h6b == _myNewVec_95_T_3[6:0] ? myVec_107 : _GEN_4372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4374 = 7'h6c == _myNewVec_95_T_3[6:0] ? myVec_108 : _GEN_4373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4375 = 7'h6d == _myNewVec_95_T_3[6:0] ? myVec_109 : _GEN_4374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4376 = 7'h6e == _myNewVec_95_T_3[6:0] ? myVec_110 : _GEN_4375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4377 = 7'h6f == _myNewVec_95_T_3[6:0] ? myVec_111 : _GEN_4376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4378 = 7'h70 == _myNewVec_95_T_3[6:0] ? myVec_112 : _GEN_4377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4379 = 7'h71 == _myNewVec_95_T_3[6:0] ? myVec_113 : _GEN_4378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4380 = 7'h72 == _myNewVec_95_T_3[6:0] ? myVec_114 : _GEN_4379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4381 = 7'h73 == _myNewVec_95_T_3[6:0] ? myVec_115 : _GEN_4380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4382 = 7'h74 == _myNewVec_95_T_3[6:0] ? myVec_116 : _GEN_4381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4383 = 7'h75 == _myNewVec_95_T_3[6:0] ? myVec_117 : _GEN_4382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4384 = 7'h76 == _myNewVec_95_T_3[6:0] ? myVec_118 : _GEN_4383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4385 = 7'h77 == _myNewVec_95_T_3[6:0] ? myVec_119 : _GEN_4384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4386 = 7'h78 == _myNewVec_95_T_3[6:0] ? myVec_120 : _GEN_4385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4387 = 7'h79 == _myNewVec_95_T_3[6:0] ? myVec_121 : _GEN_4386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4388 = 7'h7a == _myNewVec_95_T_3[6:0] ? myVec_122 : _GEN_4387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4389 = 7'h7b == _myNewVec_95_T_3[6:0] ? myVec_123 : _GEN_4388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4390 = 7'h7c == _myNewVec_95_T_3[6:0] ? myVec_124 : _GEN_4389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4391 = 7'h7d == _myNewVec_95_T_3[6:0] ? myVec_125 : _GEN_4390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4392 = 7'h7e == _myNewVec_95_T_3[6:0] ? myVec_126 : _GEN_4391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_95 = 7'h7f == _myNewVec_95_T_3[6:0] ? myVec_127 : _GEN_4392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_94_T_3 = _myNewVec_127_T_1 + 16'h21; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_4395 = 7'h1 == _myNewVec_94_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4396 = 7'h2 == _myNewVec_94_T_3[6:0] ? myVec_2 : _GEN_4395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4397 = 7'h3 == _myNewVec_94_T_3[6:0] ? myVec_3 : _GEN_4396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4398 = 7'h4 == _myNewVec_94_T_3[6:0] ? myVec_4 : _GEN_4397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4399 = 7'h5 == _myNewVec_94_T_3[6:0] ? myVec_5 : _GEN_4398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4400 = 7'h6 == _myNewVec_94_T_3[6:0] ? myVec_6 : _GEN_4399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4401 = 7'h7 == _myNewVec_94_T_3[6:0] ? myVec_7 : _GEN_4400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4402 = 7'h8 == _myNewVec_94_T_3[6:0] ? myVec_8 : _GEN_4401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4403 = 7'h9 == _myNewVec_94_T_3[6:0] ? myVec_9 : _GEN_4402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4404 = 7'ha == _myNewVec_94_T_3[6:0] ? myVec_10 : _GEN_4403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4405 = 7'hb == _myNewVec_94_T_3[6:0] ? myVec_11 : _GEN_4404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4406 = 7'hc == _myNewVec_94_T_3[6:0] ? myVec_12 : _GEN_4405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4407 = 7'hd == _myNewVec_94_T_3[6:0] ? myVec_13 : _GEN_4406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4408 = 7'he == _myNewVec_94_T_3[6:0] ? myVec_14 : _GEN_4407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4409 = 7'hf == _myNewVec_94_T_3[6:0] ? myVec_15 : _GEN_4408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4410 = 7'h10 == _myNewVec_94_T_3[6:0] ? myVec_16 : _GEN_4409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4411 = 7'h11 == _myNewVec_94_T_3[6:0] ? myVec_17 : _GEN_4410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4412 = 7'h12 == _myNewVec_94_T_3[6:0] ? myVec_18 : _GEN_4411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4413 = 7'h13 == _myNewVec_94_T_3[6:0] ? myVec_19 : _GEN_4412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4414 = 7'h14 == _myNewVec_94_T_3[6:0] ? myVec_20 : _GEN_4413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4415 = 7'h15 == _myNewVec_94_T_3[6:0] ? myVec_21 : _GEN_4414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4416 = 7'h16 == _myNewVec_94_T_3[6:0] ? myVec_22 : _GEN_4415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4417 = 7'h17 == _myNewVec_94_T_3[6:0] ? myVec_23 : _GEN_4416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4418 = 7'h18 == _myNewVec_94_T_3[6:0] ? myVec_24 : _GEN_4417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4419 = 7'h19 == _myNewVec_94_T_3[6:0] ? myVec_25 : _GEN_4418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4420 = 7'h1a == _myNewVec_94_T_3[6:0] ? myVec_26 : _GEN_4419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4421 = 7'h1b == _myNewVec_94_T_3[6:0] ? myVec_27 : _GEN_4420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4422 = 7'h1c == _myNewVec_94_T_3[6:0] ? myVec_28 : _GEN_4421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4423 = 7'h1d == _myNewVec_94_T_3[6:0] ? myVec_29 : _GEN_4422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4424 = 7'h1e == _myNewVec_94_T_3[6:0] ? myVec_30 : _GEN_4423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4425 = 7'h1f == _myNewVec_94_T_3[6:0] ? myVec_31 : _GEN_4424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4426 = 7'h20 == _myNewVec_94_T_3[6:0] ? myVec_32 : _GEN_4425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4427 = 7'h21 == _myNewVec_94_T_3[6:0] ? myVec_33 : _GEN_4426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4428 = 7'h22 == _myNewVec_94_T_3[6:0] ? myVec_34 : _GEN_4427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4429 = 7'h23 == _myNewVec_94_T_3[6:0] ? myVec_35 : _GEN_4428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4430 = 7'h24 == _myNewVec_94_T_3[6:0] ? myVec_36 : _GEN_4429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4431 = 7'h25 == _myNewVec_94_T_3[6:0] ? myVec_37 : _GEN_4430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4432 = 7'h26 == _myNewVec_94_T_3[6:0] ? myVec_38 : _GEN_4431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4433 = 7'h27 == _myNewVec_94_T_3[6:0] ? myVec_39 : _GEN_4432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4434 = 7'h28 == _myNewVec_94_T_3[6:0] ? myVec_40 : _GEN_4433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4435 = 7'h29 == _myNewVec_94_T_3[6:0] ? myVec_41 : _GEN_4434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4436 = 7'h2a == _myNewVec_94_T_3[6:0] ? myVec_42 : _GEN_4435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4437 = 7'h2b == _myNewVec_94_T_3[6:0] ? myVec_43 : _GEN_4436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4438 = 7'h2c == _myNewVec_94_T_3[6:0] ? myVec_44 : _GEN_4437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4439 = 7'h2d == _myNewVec_94_T_3[6:0] ? myVec_45 : _GEN_4438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4440 = 7'h2e == _myNewVec_94_T_3[6:0] ? myVec_46 : _GEN_4439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4441 = 7'h2f == _myNewVec_94_T_3[6:0] ? myVec_47 : _GEN_4440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4442 = 7'h30 == _myNewVec_94_T_3[6:0] ? myVec_48 : _GEN_4441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4443 = 7'h31 == _myNewVec_94_T_3[6:0] ? myVec_49 : _GEN_4442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4444 = 7'h32 == _myNewVec_94_T_3[6:0] ? myVec_50 : _GEN_4443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4445 = 7'h33 == _myNewVec_94_T_3[6:0] ? myVec_51 : _GEN_4444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4446 = 7'h34 == _myNewVec_94_T_3[6:0] ? myVec_52 : _GEN_4445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4447 = 7'h35 == _myNewVec_94_T_3[6:0] ? myVec_53 : _GEN_4446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4448 = 7'h36 == _myNewVec_94_T_3[6:0] ? myVec_54 : _GEN_4447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4449 = 7'h37 == _myNewVec_94_T_3[6:0] ? myVec_55 : _GEN_4448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4450 = 7'h38 == _myNewVec_94_T_3[6:0] ? myVec_56 : _GEN_4449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4451 = 7'h39 == _myNewVec_94_T_3[6:0] ? myVec_57 : _GEN_4450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4452 = 7'h3a == _myNewVec_94_T_3[6:0] ? myVec_58 : _GEN_4451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4453 = 7'h3b == _myNewVec_94_T_3[6:0] ? myVec_59 : _GEN_4452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4454 = 7'h3c == _myNewVec_94_T_3[6:0] ? myVec_60 : _GEN_4453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4455 = 7'h3d == _myNewVec_94_T_3[6:0] ? myVec_61 : _GEN_4454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4456 = 7'h3e == _myNewVec_94_T_3[6:0] ? myVec_62 : _GEN_4455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4457 = 7'h3f == _myNewVec_94_T_3[6:0] ? myVec_63 : _GEN_4456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4458 = 7'h40 == _myNewVec_94_T_3[6:0] ? myVec_64 : _GEN_4457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4459 = 7'h41 == _myNewVec_94_T_3[6:0] ? myVec_65 : _GEN_4458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4460 = 7'h42 == _myNewVec_94_T_3[6:0] ? myVec_66 : _GEN_4459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4461 = 7'h43 == _myNewVec_94_T_3[6:0] ? myVec_67 : _GEN_4460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4462 = 7'h44 == _myNewVec_94_T_3[6:0] ? myVec_68 : _GEN_4461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4463 = 7'h45 == _myNewVec_94_T_3[6:0] ? myVec_69 : _GEN_4462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4464 = 7'h46 == _myNewVec_94_T_3[6:0] ? myVec_70 : _GEN_4463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4465 = 7'h47 == _myNewVec_94_T_3[6:0] ? myVec_71 : _GEN_4464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4466 = 7'h48 == _myNewVec_94_T_3[6:0] ? myVec_72 : _GEN_4465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4467 = 7'h49 == _myNewVec_94_T_3[6:0] ? myVec_73 : _GEN_4466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4468 = 7'h4a == _myNewVec_94_T_3[6:0] ? myVec_74 : _GEN_4467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4469 = 7'h4b == _myNewVec_94_T_3[6:0] ? myVec_75 : _GEN_4468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4470 = 7'h4c == _myNewVec_94_T_3[6:0] ? myVec_76 : _GEN_4469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4471 = 7'h4d == _myNewVec_94_T_3[6:0] ? myVec_77 : _GEN_4470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4472 = 7'h4e == _myNewVec_94_T_3[6:0] ? myVec_78 : _GEN_4471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4473 = 7'h4f == _myNewVec_94_T_3[6:0] ? myVec_79 : _GEN_4472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4474 = 7'h50 == _myNewVec_94_T_3[6:0] ? myVec_80 : _GEN_4473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4475 = 7'h51 == _myNewVec_94_T_3[6:0] ? myVec_81 : _GEN_4474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4476 = 7'h52 == _myNewVec_94_T_3[6:0] ? myVec_82 : _GEN_4475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4477 = 7'h53 == _myNewVec_94_T_3[6:0] ? myVec_83 : _GEN_4476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4478 = 7'h54 == _myNewVec_94_T_3[6:0] ? myVec_84 : _GEN_4477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4479 = 7'h55 == _myNewVec_94_T_3[6:0] ? myVec_85 : _GEN_4478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4480 = 7'h56 == _myNewVec_94_T_3[6:0] ? myVec_86 : _GEN_4479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4481 = 7'h57 == _myNewVec_94_T_3[6:0] ? myVec_87 : _GEN_4480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4482 = 7'h58 == _myNewVec_94_T_3[6:0] ? myVec_88 : _GEN_4481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4483 = 7'h59 == _myNewVec_94_T_3[6:0] ? myVec_89 : _GEN_4482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4484 = 7'h5a == _myNewVec_94_T_3[6:0] ? myVec_90 : _GEN_4483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4485 = 7'h5b == _myNewVec_94_T_3[6:0] ? myVec_91 : _GEN_4484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4486 = 7'h5c == _myNewVec_94_T_3[6:0] ? myVec_92 : _GEN_4485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4487 = 7'h5d == _myNewVec_94_T_3[6:0] ? myVec_93 : _GEN_4486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4488 = 7'h5e == _myNewVec_94_T_3[6:0] ? myVec_94 : _GEN_4487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4489 = 7'h5f == _myNewVec_94_T_3[6:0] ? myVec_95 : _GEN_4488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4490 = 7'h60 == _myNewVec_94_T_3[6:0] ? myVec_96 : _GEN_4489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4491 = 7'h61 == _myNewVec_94_T_3[6:0] ? myVec_97 : _GEN_4490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4492 = 7'h62 == _myNewVec_94_T_3[6:0] ? myVec_98 : _GEN_4491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4493 = 7'h63 == _myNewVec_94_T_3[6:0] ? myVec_99 : _GEN_4492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4494 = 7'h64 == _myNewVec_94_T_3[6:0] ? myVec_100 : _GEN_4493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4495 = 7'h65 == _myNewVec_94_T_3[6:0] ? myVec_101 : _GEN_4494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4496 = 7'h66 == _myNewVec_94_T_3[6:0] ? myVec_102 : _GEN_4495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4497 = 7'h67 == _myNewVec_94_T_3[6:0] ? myVec_103 : _GEN_4496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4498 = 7'h68 == _myNewVec_94_T_3[6:0] ? myVec_104 : _GEN_4497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4499 = 7'h69 == _myNewVec_94_T_3[6:0] ? myVec_105 : _GEN_4498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4500 = 7'h6a == _myNewVec_94_T_3[6:0] ? myVec_106 : _GEN_4499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4501 = 7'h6b == _myNewVec_94_T_3[6:0] ? myVec_107 : _GEN_4500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4502 = 7'h6c == _myNewVec_94_T_3[6:0] ? myVec_108 : _GEN_4501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4503 = 7'h6d == _myNewVec_94_T_3[6:0] ? myVec_109 : _GEN_4502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4504 = 7'h6e == _myNewVec_94_T_3[6:0] ? myVec_110 : _GEN_4503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4505 = 7'h6f == _myNewVec_94_T_3[6:0] ? myVec_111 : _GEN_4504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4506 = 7'h70 == _myNewVec_94_T_3[6:0] ? myVec_112 : _GEN_4505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4507 = 7'h71 == _myNewVec_94_T_3[6:0] ? myVec_113 : _GEN_4506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4508 = 7'h72 == _myNewVec_94_T_3[6:0] ? myVec_114 : _GEN_4507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4509 = 7'h73 == _myNewVec_94_T_3[6:0] ? myVec_115 : _GEN_4508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4510 = 7'h74 == _myNewVec_94_T_3[6:0] ? myVec_116 : _GEN_4509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4511 = 7'h75 == _myNewVec_94_T_3[6:0] ? myVec_117 : _GEN_4510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4512 = 7'h76 == _myNewVec_94_T_3[6:0] ? myVec_118 : _GEN_4511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4513 = 7'h77 == _myNewVec_94_T_3[6:0] ? myVec_119 : _GEN_4512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4514 = 7'h78 == _myNewVec_94_T_3[6:0] ? myVec_120 : _GEN_4513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4515 = 7'h79 == _myNewVec_94_T_3[6:0] ? myVec_121 : _GEN_4514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4516 = 7'h7a == _myNewVec_94_T_3[6:0] ? myVec_122 : _GEN_4515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4517 = 7'h7b == _myNewVec_94_T_3[6:0] ? myVec_123 : _GEN_4516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4518 = 7'h7c == _myNewVec_94_T_3[6:0] ? myVec_124 : _GEN_4517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4519 = 7'h7d == _myNewVec_94_T_3[6:0] ? myVec_125 : _GEN_4518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4520 = 7'h7e == _myNewVec_94_T_3[6:0] ? myVec_126 : _GEN_4519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_94 = 7'h7f == _myNewVec_94_T_3[6:0] ? myVec_127 : _GEN_4520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_93_T_3 = _myNewVec_127_T_1 + 16'h22; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_4523 = 7'h1 == _myNewVec_93_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4524 = 7'h2 == _myNewVec_93_T_3[6:0] ? myVec_2 : _GEN_4523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4525 = 7'h3 == _myNewVec_93_T_3[6:0] ? myVec_3 : _GEN_4524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4526 = 7'h4 == _myNewVec_93_T_3[6:0] ? myVec_4 : _GEN_4525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4527 = 7'h5 == _myNewVec_93_T_3[6:0] ? myVec_5 : _GEN_4526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4528 = 7'h6 == _myNewVec_93_T_3[6:0] ? myVec_6 : _GEN_4527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4529 = 7'h7 == _myNewVec_93_T_3[6:0] ? myVec_7 : _GEN_4528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4530 = 7'h8 == _myNewVec_93_T_3[6:0] ? myVec_8 : _GEN_4529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4531 = 7'h9 == _myNewVec_93_T_3[6:0] ? myVec_9 : _GEN_4530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4532 = 7'ha == _myNewVec_93_T_3[6:0] ? myVec_10 : _GEN_4531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4533 = 7'hb == _myNewVec_93_T_3[6:0] ? myVec_11 : _GEN_4532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4534 = 7'hc == _myNewVec_93_T_3[6:0] ? myVec_12 : _GEN_4533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4535 = 7'hd == _myNewVec_93_T_3[6:0] ? myVec_13 : _GEN_4534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4536 = 7'he == _myNewVec_93_T_3[6:0] ? myVec_14 : _GEN_4535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4537 = 7'hf == _myNewVec_93_T_3[6:0] ? myVec_15 : _GEN_4536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4538 = 7'h10 == _myNewVec_93_T_3[6:0] ? myVec_16 : _GEN_4537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4539 = 7'h11 == _myNewVec_93_T_3[6:0] ? myVec_17 : _GEN_4538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4540 = 7'h12 == _myNewVec_93_T_3[6:0] ? myVec_18 : _GEN_4539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4541 = 7'h13 == _myNewVec_93_T_3[6:0] ? myVec_19 : _GEN_4540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4542 = 7'h14 == _myNewVec_93_T_3[6:0] ? myVec_20 : _GEN_4541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4543 = 7'h15 == _myNewVec_93_T_3[6:0] ? myVec_21 : _GEN_4542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4544 = 7'h16 == _myNewVec_93_T_3[6:0] ? myVec_22 : _GEN_4543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4545 = 7'h17 == _myNewVec_93_T_3[6:0] ? myVec_23 : _GEN_4544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4546 = 7'h18 == _myNewVec_93_T_3[6:0] ? myVec_24 : _GEN_4545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4547 = 7'h19 == _myNewVec_93_T_3[6:0] ? myVec_25 : _GEN_4546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4548 = 7'h1a == _myNewVec_93_T_3[6:0] ? myVec_26 : _GEN_4547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4549 = 7'h1b == _myNewVec_93_T_3[6:0] ? myVec_27 : _GEN_4548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4550 = 7'h1c == _myNewVec_93_T_3[6:0] ? myVec_28 : _GEN_4549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4551 = 7'h1d == _myNewVec_93_T_3[6:0] ? myVec_29 : _GEN_4550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4552 = 7'h1e == _myNewVec_93_T_3[6:0] ? myVec_30 : _GEN_4551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4553 = 7'h1f == _myNewVec_93_T_3[6:0] ? myVec_31 : _GEN_4552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4554 = 7'h20 == _myNewVec_93_T_3[6:0] ? myVec_32 : _GEN_4553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4555 = 7'h21 == _myNewVec_93_T_3[6:0] ? myVec_33 : _GEN_4554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4556 = 7'h22 == _myNewVec_93_T_3[6:0] ? myVec_34 : _GEN_4555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4557 = 7'h23 == _myNewVec_93_T_3[6:0] ? myVec_35 : _GEN_4556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4558 = 7'h24 == _myNewVec_93_T_3[6:0] ? myVec_36 : _GEN_4557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4559 = 7'h25 == _myNewVec_93_T_3[6:0] ? myVec_37 : _GEN_4558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4560 = 7'h26 == _myNewVec_93_T_3[6:0] ? myVec_38 : _GEN_4559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4561 = 7'h27 == _myNewVec_93_T_3[6:0] ? myVec_39 : _GEN_4560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4562 = 7'h28 == _myNewVec_93_T_3[6:0] ? myVec_40 : _GEN_4561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4563 = 7'h29 == _myNewVec_93_T_3[6:0] ? myVec_41 : _GEN_4562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4564 = 7'h2a == _myNewVec_93_T_3[6:0] ? myVec_42 : _GEN_4563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4565 = 7'h2b == _myNewVec_93_T_3[6:0] ? myVec_43 : _GEN_4564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4566 = 7'h2c == _myNewVec_93_T_3[6:0] ? myVec_44 : _GEN_4565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4567 = 7'h2d == _myNewVec_93_T_3[6:0] ? myVec_45 : _GEN_4566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4568 = 7'h2e == _myNewVec_93_T_3[6:0] ? myVec_46 : _GEN_4567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4569 = 7'h2f == _myNewVec_93_T_3[6:0] ? myVec_47 : _GEN_4568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4570 = 7'h30 == _myNewVec_93_T_3[6:0] ? myVec_48 : _GEN_4569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4571 = 7'h31 == _myNewVec_93_T_3[6:0] ? myVec_49 : _GEN_4570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4572 = 7'h32 == _myNewVec_93_T_3[6:0] ? myVec_50 : _GEN_4571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4573 = 7'h33 == _myNewVec_93_T_3[6:0] ? myVec_51 : _GEN_4572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4574 = 7'h34 == _myNewVec_93_T_3[6:0] ? myVec_52 : _GEN_4573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4575 = 7'h35 == _myNewVec_93_T_3[6:0] ? myVec_53 : _GEN_4574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4576 = 7'h36 == _myNewVec_93_T_3[6:0] ? myVec_54 : _GEN_4575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4577 = 7'h37 == _myNewVec_93_T_3[6:0] ? myVec_55 : _GEN_4576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4578 = 7'h38 == _myNewVec_93_T_3[6:0] ? myVec_56 : _GEN_4577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4579 = 7'h39 == _myNewVec_93_T_3[6:0] ? myVec_57 : _GEN_4578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4580 = 7'h3a == _myNewVec_93_T_3[6:0] ? myVec_58 : _GEN_4579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4581 = 7'h3b == _myNewVec_93_T_3[6:0] ? myVec_59 : _GEN_4580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4582 = 7'h3c == _myNewVec_93_T_3[6:0] ? myVec_60 : _GEN_4581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4583 = 7'h3d == _myNewVec_93_T_3[6:0] ? myVec_61 : _GEN_4582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4584 = 7'h3e == _myNewVec_93_T_3[6:0] ? myVec_62 : _GEN_4583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4585 = 7'h3f == _myNewVec_93_T_3[6:0] ? myVec_63 : _GEN_4584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4586 = 7'h40 == _myNewVec_93_T_3[6:0] ? myVec_64 : _GEN_4585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4587 = 7'h41 == _myNewVec_93_T_3[6:0] ? myVec_65 : _GEN_4586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4588 = 7'h42 == _myNewVec_93_T_3[6:0] ? myVec_66 : _GEN_4587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4589 = 7'h43 == _myNewVec_93_T_3[6:0] ? myVec_67 : _GEN_4588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4590 = 7'h44 == _myNewVec_93_T_3[6:0] ? myVec_68 : _GEN_4589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4591 = 7'h45 == _myNewVec_93_T_3[6:0] ? myVec_69 : _GEN_4590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4592 = 7'h46 == _myNewVec_93_T_3[6:0] ? myVec_70 : _GEN_4591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4593 = 7'h47 == _myNewVec_93_T_3[6:0] ? myVec_71 : _GEN_4592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4594 = 7'h48 == _myNewVec_93_T_3[6:0] ? myVec_72 : _GEN_4593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4595 = 7'h49 == _myNewVec_93_T_3[6:0] ? myVec_73 : _GEN_4594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4596 = 7'h4a == _myNewVec_93_T_3[6:0] ? myVec_74 : _GEN_4595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4597 = 7'h4b == _myNewVec_93_T_3[6:0] ? myVec_75 : _GEN_4596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4598 = 7'h4c == _myNewVec_93_T_3[6:0] ? myVec_76 : _GEN_4597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4599 = 7'h4d == _myNewVec_93_T_3[6:0] ? myVec_77 : _GEN_4598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4600 = 7'h4e == _myNewVec_93_T_3[6:0] ? myVec_78 : _GEN_4599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4601 = 7'h4f == _myNewVec_93_T_3[6:0] ? myVec_79 : _GEN_4600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4602 = 7'h50 == _myNewVec_93_T_3[6:0] ? myVec_80 : _GEN_4601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4603 = 7'h51 == _myNewVec_93_T_3[6:0] ? myVec_81 : _GEN_4602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4604 = 7'h52 == _myNewVec_93_T_3[6:0] ? myVec_82 : _GEN_4603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4605 = 7'h53 == _myNewVec_93_T_3[6:0] ? myVec_83 : _GEN_4604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4606 = 7'h54 == _myNewVec_93_T_3[6:0] ? myVec_84 : _GEN_4605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4607 = 7'h55 == _myNewVec_93_T_3[6:0] ? myVec_85 : _GEN_4606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4608 = 7'h56 == _myNewVec_93_T_3[6:0] ? myVec_86 : _GEN_4607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4609 = 7'h57 == _myNewVec_93_T_3[6:0] ? myVec_87 : _GEN_4608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4610 = 7'h58 == _myNewVec_93_T_3[6:0] ? myVec_88 : _GEN_4609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4611 = 7'h59 == _myNewVec_93_T_3[6:0] ? myVec_89 : _GEN_4610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4612 = 7'h5a == _myNewVec_93_T_3[6:0] ? myVec_90 : _GEN_4611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4613 = 7'h5b == _myNewVec_93_T_3[6:0] ? myVec_91 : _GEN_4612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4614 = 7'h5c == _myNewVec_93_T_3[6:0] ? myVec_92 : _GEN_4613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4615 = 7'h5d == _myNewVec_93_T_3[6:0] ? myVec_93 : _GEN_4614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4616 = 7'h5e == _myNewVec_93_T_3[6:0] ? myVec_94 : _GEN_4615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4617 = 7'h5f == _myNewVec_93_T_3[6:0] ? myVec_95 : _GEN_4616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4618 = 7'h60 == _myNewVec_93_T_3[6:0] ? myVec_96 : _GEN_4617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4619 = 7'h61 == _myNewVec_93_T_3[6:0] ? myVec_97 : _GEN_4618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4620 = 7'h62 == _myNewVec_93_T_3[6:0] ? myVec_98 : _GEN_4619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4621 = 7'h63 == _myNewVec_93_T_3[6:0] ? myVec_99 : _GEN_4620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4622 = 7'h64 == _myNewVec_93_T_3[6:0] ? myVec_100 : _GEN_4621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4623 = 7'h65 == _myNewVec_93_T_3[6:0] ? myVec_101 : _GEN_4622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4624 = 7'h66 == _myNewVec_93_T_3[6:0] ? myVec_102 : _GEN_4623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4625 = 7'h67 == _myNewVec_93_T_3[6:0] ? myVec_103 : _GEN_4624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4626 = 7'h68 == _myNewVec_93_T_3[6:0] ? myVec_104 : _GEN_4625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4627 = 7'h69 == _myNewVec_93_T_3[6:0] ? myVec_105 : _GEN_4626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4628 = 7'h6a == _myNewVec_93_T_3[6:0] ? myVec_106 : _GEN_4627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4629 = 7'h6b == _myNewVec_93_T_3[6:0] ? myVec_107 : _GEN_4628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4630 = 7'h6c == _myNewVec_93_T_3[6:0] ? myVec_108 : _GEN_4629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4631 = 7'h6d == _myNewVec_93_T_3[6:0] ? myVec_109 : _GEN_4630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4632 = 7'h6e == _myNewVec_93_T_3[6:0] ? myVec_110 : _GEN_4631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4633 = 7'h6f == _myNewVec_93_T_3[6:0] ? myVec_111 : _GEN_4632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4634 = 7'h70 == _myNewVec_93_T_3[6:0] ? myVec_112 : _GEN_4633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4635 = 7'h71 == _myNewVec_93_T_3[6:0] ? myVec_113 : _GEN_4634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4636 = 7'h72 == _myNewVec_93_T_3[6:0] ? myVec_114 : _GEN_4635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4637 = 7'h73 == _myNewVec_93_T_3[6:0] ? myVec_115 : _GEN_4636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4638 = 7'h74 == _myNewVec_93_T_3[6:0] ? myVec_116 : _GEN_4637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4639 = 7'h75 == _myNewVec_93_T_3[6:0] ? myVec_117 : _GEN_4638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4640 = 7'h76 == _myNewVec_93_T_3[6:0] ? myVec_118 : _GEN_4639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4641 = 7'h77 == _myNewVec_93_T_3[6:0] ? myVec_119 : _GEN_4640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4642 = 7'h78 == _myNewVec_93_T_3[6:0] ? myVec_120 : _GEN_4641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4643 = 7'h79 == _myNewVec_93_T_3[6:0] ? myVec_121 : _GEN_4642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4644 = 7'h7a == _myNewVec_93_T_3[6:0] ? myVec_122 : _GEN_4643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4645 = 7'h7b == _myNewVec_93_T_3[6:0] ? myVec_123 : _GEN_4644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4646 = 7'h7c == _myNewVec_93_T_3[6:0] ? myVec_124 : _GEN_4645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4647 = 7'h7d == _myNewVec_93_T_3[6:0] ? myVec_125 : _GEN_4646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4648 = 7'h7e == _myNewVec_93_T_3[6:0] ? myVec_126 : _GEN_4647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_93 = 7'h7f == _myNewVec_93_T_3[6:0] ? myVec_127 : _GEN_4648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_92_T_3 = _myNewVec_127_T_1 + 16'h23; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_4651 = 7'h1 == _myNewVec_92_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4652 = 7'h2 == _myNewVec_92_T_3[6:0] ? myVec_2 : _GEN_4651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4653 = 7'h3 == _myNewVec_92_T_3[6:0] ? myVec_3 : _GEN_4652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4654 = 7'h4 == _myNewVec_92_T_3[6:0] ? myVec_4 : _GEN_4653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4655 = 7'h5 == _myNewVec_92_T_3[6:0] ? myVec_5 : _GEN_4654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4656 = 7'h6 == _myNewVec_92_T_3[6:0] ? myVec_6 : _GEN_4655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4657 = 7'h7 == _myNewVec_92_T_3[6:0] ? myVec_7 : _GEN_4656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4658 = 7'h8 == _myNewVec_92_T_3[6:0] ? myVec_8 : _GEN_4657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4659 = 7'h9 == _myNewVec_92_T_3[6:0] ? myVec_9 : _GEN_4658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4660 = 7'ha == _myNewVec_92_T_3[6:0] ? myVec_10 : _GEN_4659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4661 = 7'hb == _myNewVec_92_T_3[6:0] ? myVec_11 : _GEN_4660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4662 = 7'hc == _myNewVec_92_T_3[6:0] ? myVec_12 : _GEN_4661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4663 = 7'hd == _myNewVec_92_T_3[6:0] ? myVec_13 : _GEN_4662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4664 = 7'he == _myNewVec_92_T_3[6:0] ? myVec_14 : _GEN_4663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4665 = 7'hf == _myNewVec_92_T_3[6:0] ? myVec_15 : _GEN_4664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4666 = 7'h10 == _myNewVec_92_T_3[6:0] ? myVec_16 : _GEN_4665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4667 = 7'h11 == _myNewVec_92_T_3[6:0] ? myVec_17 : _GEN_4666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4668 = 7'h12 == _myNewVec_92_T_3[6:0] ? myVec_18 : _GEN_4667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4669 = 7'h13 == _myNewVec_92_T_3[6:0] ? myVec_19 : _GEN_4668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4670 = 7'h14 == _myNewVec_92_T_3[6:0] ? myVec_20 : _GEN_4669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4671 = 7'h15 == _myNewVec_92_T_3[6:0] ? myVec_21 : _GEN_4670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4672 = 7'h16 == _myNewVec_92_T_3[6:0] ? myVec_22 : _GEN_4671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4673 = 7'h17 == _myNewVec_92_T_3[6:0] ? myVec_23 : _GEN_4672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4674 = 7'h18 == _myNewVec_92_T_3[6:0] ? myVec_24 : _GEN_4673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4675 = 7'h19 == _myNewVec_92_T_3[6:0] ? myVec_25 : _GEN_4674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4676 = 7'h1a == _myNewVec_92_T_3[6:0] ? myVec_26 : _GEN_4675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4677 = 7'h1b == _myNewVec_92_T_3[6:0] ? myVec_27 : _GEN_4676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4678 = 7'h1c == _myNewVec_92_T_3[6:0] ? myVec_28 : _GEN_4677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4679 = 7'h1d == _myNewVec_92_T_3[6:0] ? myVec_29 : _GEN_4678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4680 = 7'h1e == _myNewVec_92_T_3[6:0] ? myVec_30 : _GEN_4679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4681 = 7'h1f == _myNewVec_92_T_3[6:0] ? myVec_31 : _GEN_4680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4682 = 7'h20 == _myNewVec_92_T_3[6:0] ? myVec_32 : _GEN_4681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4683 = 7'h21 == _myNewVec_92_T_3[6:0] ? myVec_33 : _GEN_4682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4684 = 7'h22 == _myNewVec_92_T_3[6:0] ? myVec_34 : _GEN_4683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4685 = 7'h23 == _myNewVec_92_T_3[6:0] ? myVec_35 : _GEN_4684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4686 = 7'h24 == _myNewVec_92_T_3[6:0] ? myVec_36 : _GEN_4685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4687 = 7'h25 == _myNewVec_92_T_3[6:0] ? myVec_37 : _GEN_4686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4688 = 7'h26 == _myNewVec_92_T_3[6:0] ? myVec_38 : _GEN_4687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4689 = 7'h27 == _myNewVec_92_T_3[6:0] ? myVec_39 : _GEN_4688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4690 = 7'h28 == _myNewVec_92_T_3[6:0] ? myVec_40 : _GEN_4689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4691 = 7'h29 == _myNewVec_92_T_3[6:0] ? myVec_41 : _GEN_4690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4692 = 7'h2a == _myNewVec_92_T_3[6:0] ? myVec_42 : _GEN_4691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4693 = 7'h2b == _myNewVec_92_T_3[6:0] ? myVec_43 : _GEN_4692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4694 = 7'h2c == _myNewVec_92_T_3[6:0] ? myVec_44 : _GEN_4693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4695 = 7'h2d == _myNewVec_92_T_3[6:0] ? myVec_45 : _GEN_4694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4696 = 7'h2e == _myNewVec_92_T_3[6:0] ? myVec_46 : _GEN_4695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4697 = 7'h2f == _myNewVec_92_T_3[6:0] ? myVec_47 : _GEN_4696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4698 = 7'h30 == _myNewVec_92_T_3[6:0] ? myVec_48 : _GEN_4697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4699 = 7'h31 == _myNewVec_92_T_3[6:0] ? myVec_49 : _GEN_4698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4700 = 7'h32 == _myNewVec_92_T_3[6:0] ? myVec_50 : _GEN_4699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4701 = 7'h33 == _myNewVec_92_T_3[6:0] ? myVec_51 : _GEN_4700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4702 = 7'h34 == _myNewVec_92_T_3[6:0] ? myVec_52 : _GEN_4701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4703 = 7'h35 == _myNewVec_92_T_3[6:0] ? myVec_53 : _GEN_4702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4704 = 7'h36 == _myNewVec_92_T_3[6:0] ? myVec_54 : _GEN_4703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4705 = 7'h37 == _myNewVec_92_T_3[6:0] ? myVec_55 : _GEN_4704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4706 = 7'h38 == _myNewVec_92_T_3[6:0] ? myVec_56 : _GEN_4705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4707 = 7'h39 == _myNewVec_92_T_3[6:0] ? myVec_57 : _GEN_4706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4708 = 7'h3a == _myNewVec_92_T_3[6:0] ? myVec_58 : _GEN_4707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4709 = 7'h3b == _myNewVec_92_T_3[6:0] ? myVec_59 : _GEN_4708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4710 = 7'h3c == _myNewVec_92_T_3[6:0] ? myVec_60 : _GEN_4709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4711 = 7'h3d == _myNewVec_92_T_3[6:0] ? myVec_61 : _GEN_4710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4712 = 7'h3e == _myNewVec_92_T_3[6:0] ? myVec_62 : _GEN_4711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4713 = 7'h3f == _myNewVec_92_T_3[6:0] ? myVec_63 : _GEN_4712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4714 = 7'h40 == _myNewVec_92_T_3[6:0] ? myVec_64 : _GEN_4713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4715 = 7'h41 == _myNewVec_92_T_3[6:0] ? myVec_65 : _GEN_4714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4716 = 7'h42 == _myNewVec_92_T_3[6:0] ? myVec_66 : _GEN_4715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4717 = 7'h43 == _myNewVec_92_T_3[6:0] ? myVec_67 : _GEN_4716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4718 = 7'h44 == _myNewVec_92_T_3[6:0] ? myVec_68 : _GEN_4717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4719 = 7'h45 == _myNewVec_92_T_3[6:0] ? myVec_69 : _GEN_4718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4720 = 7'h46 == _myNewVec_92_T_3[6:0] ? myVec_70 : _GEN_4719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4721 = 7'h47 == _myNewVec_92_T_3[6:0] ? myVec_71 : _GEN_4720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4722 = 7'h48 == _myNewVec_92_T_3[6:0] ? myVec_72 : _GEN_4721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4723 = 7'h49 == _myNewVec_92_T_3[6:0] ? myVec_73 : _GEN_4722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4724 = 7'h4a == _myNewVec_92_T_3[6:0] ? myVec_74 : _GEN_4723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4725 = 7'h4b == _myNewVec_92_T_3[6:0] ? myVec_75 : _GEN_4724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4726 = 7'h4c == _myNewVec_92_T_3[6:0] ? myVec_76 : _GEN_4725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4727 = 7'h4d == _myNewVec_92_T_3[6:0] ? myVec_77 : _GEN_4726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4728 = 7'h4e == _myNewVec_92_T_3[6:0] ? myVec_78 : _GEN_4727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4729 = 7'h4f == _myNewVec_92_T_3[6:0] ? myVec_79 : _GEN_4728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4730 = 7'h50 == _myNewVec_92_T_3[6:0] ? myVec_80 : _GEN_4729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4731 = 7'h51 == _myNewVec_92_T_3[6:0] ? myVec_81 : _GEN_4730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4732 = 7'h52 == _myNewVec_92_T_3[6:0] ? myVec_82 : _GEN_4731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4733 = 7'h53 == _myNewVec_92_T_3[6:0] ? myVec_83 : _GEN_4732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4734 = 7'h54 == _myNewVec_92_T_3[6:0] ? myVec_84 : _GEN_4733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4735 = 7'h55 == _myNewVec_92_T_3[6:0] ? myVec_85 : _GEN_4734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4736 = 7'h56 == _myNewVec_92_T_3[6:0] ? myVec_86 : _GEN_4735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4737 = 7'h57 == _myNewVec_92_T_3[6:0] ? myVec_87 : _GEN_4736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4738 = 7'h58 == _myNewVec_92_T_3[6:0] ? myVec_88 : _GEN_4737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4739 = 7'h59 == _myNewVec_92_T_3[6:0] ? myVec_89 : _GEN_4738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4740 = 7'h5a == _myNewVec_92_T_3[6:0] ? myVec_90 : _GEN_4739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4741 = 7'h5b == _myNewVec_92_T_3[6:0] ? myVec_91 : _GEN_4740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4742 = 7'h5c == _myNewVec_92_T_3[6:0] ? myVec_92 : _GEN_4741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4743 = 7'h5d == _myNewVec_92_T_3[6:0] ? myVec_93 : _GEN_4742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4744 = 7'h5e == _myNewVec_92_T_3[6:0] ? myVec_94 : _GEN_4743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4745 = 7'h5f == _myNewVec_92_T_3[6:0] ? myVec_95 : _GEN_4744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4746 = 7'h60 == _myNewVec_92_T_3[6:0] ? myVec_96 : _GEN_4745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4747 = 7'h61 == _myNewVec_92_T_3[6:0] ? myVec_97 : _GEN_4746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4748 = 7'h62 == _myNewVec_92_T_3[6:0] ? myVec_98 : _GEN_4747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4749 = 7'h63 == _myNewVec_92_T_3[6:0] ? myVec_99 : _GEN_4748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4750 = 7'h64 == _myNewVec_92_T_3[6:0] ? myVec_100 : _GEN_4749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4751 = 7'h65 == _myNewVec_92_T_3[6:0] ? myVec_101 : _GEN_4750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4752 = 7'h66 == _myNewVec_92_T_3[6:0] ? myVec_102 : _GEN_4751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4753 = 7'h67 == _myNewVec_92_T_3[6:0] ? myVec_103 : _GEN_4752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4754 = 7'h68 == _myNewVec_92_T_3[6:0] ? myVec_104 : _GEN_4753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4755 = 7'h69 == _myNewVec_92_T_3[6:0] ? myVec_105 : _GEN_4754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4756 = 7'h6a == _myNewVec_92_T_3[6:0] ? myVec_106 : _GEN_4755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4757 = 7'h6b == _myNewVec_92_T_3[6:0] ? myVec_107 : _GEN_4756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4758 = 7'h6c == _myNewVec_92_T_3[6:0] ? myVec_108 : _GEN_4757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4759 = 7'h6d == _myNewVec_92_T_3[6:0] ? myVec_109 : _GEN_4758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4760 = 7'h6e == _myNewVec_92_T_3[6:0] ? myVec_110 : _GEN_4759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4761 = 7'h6f == _myNewVec_92_T_3[6:0] ? myVec_111 : _GEN_4760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4762 = 7'h70 == _myNewVec_92_T_3[6:0] ? myVec_112 : _GEN_4761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4763 = 7'h71 == _myNewVec_92_T_3[6:0] ? myVec_113 : _GEN_4762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4764 = 7'h72 == _myNewVec_92_T_3[6:0] ? myVec_114 : _GEN_4763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4765 = 7'h73 == _myNewVec_92_T_3[6:0] ? myVec_115 : _GEN_4764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4766 = 7'h74 == _myNewVec_92_T_3[6:0] ? myVec_116 : _GEN_4765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4767 = 7'h75 == _myNewVec_92_T_3[6:0] ? myVec_117 : _GEN_4766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4768 = 7'h76 == _myNewVec_92_T_3[6:0] ? myVec_118 : _GEN_4767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4769 = 7'h77 == _myNewVec_92_T_3[6:0] ? myVec_119 : _GEN_4768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4770 = 7'h78 == _myNewVec_92_T_3[6:0] ? myVec_120 : _GEN_4769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4771 = 7'h79 == _myNewVec_92_T_3[6:0] ? myVec_121 : _GEN_4770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4772 = 7'h7a == _myNewVec_92_T_3[6:0] ? myVec_122 : _GEN_4771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4773 = 7'h7b == _myNewVec_92_T_3[6:0] ? myVec_123 : _GEN_4772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4774 = 7'h7c == _myNewVec_92_T_3[6:0] ? myVec_124 : _GEN_4773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4775 = 7'h7d == _myNewVec_92_T_3[6:0] ? myVec_125 : _GEN_4774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4776 = 7'h7e == _myNewVec_92_T_3[6:0] ? myVec_126 : _GEN_4775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_92 = 7'h7f == _myNewVec_92_T_3[6:0] ? myVec_127 : _GEN_4776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_91_T_3 = _myNewVec_127_T_1 + 16'h24; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_4779 = 7'h1 == _myNewVec_91_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4780 = 7'h2 == _myNewVec_91_T_3[6:0] ? myVec_2 : _GEN_4779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4781 = 7'h3 == _myNewVec_91_T_3[6:0] ? myVec_3 : _GEN_4780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4782 = 7'h4 == _myNewVec_91_T_3[6:0] ? myVec_4 : _GEN_4781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4783 = 7'h5 == _myNewVec_91_T_3[6:0] ? myVec_5 : _GEN_4782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4784 = 7'h6 == _myNewVec_91_T_3[6:0] ? myVec_6 : _GEN_4783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4785 = 7'h7 == _myNewVec_91_T_3[6:0] ? myVec_7 : _GEN_4784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4786 = 7'h8 == _myNewVec_91_T_3[6:0] ? myVec_8 : _GEN_4785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4787 = 7'h9 == _myNewVec_91_T_3[6:0] ? myVec_9 : _GEN_4786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4788 = 7'ha == _myNewVec_91_T_3[6:0] ? myVec_10 : _GEN_4787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4789 = 7'hb == _myNewVec_91_T_3[6:0] ? myVec_11 : _GEN_4788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4790 = 7'hc == _myNewVec_91_T_3[6:0] ? myVec_12 : _GEN_4789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4791 = 7'hd == _myNewVec_91_T_3[6:0] ? myVec_13 : _GEN_4790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4792 = 7'he == _myNewVec_91_T_3[6:0] ? myVec_14 : _GEN_4791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4793 = 7'hf == _myNewVec_91_T_3[6:0] ? myVec_15 : _GEN_4792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4794 = 7'h10 == _myNewVec_91_T_3[6:0] ? myVec_16 : _GEN_4793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4795 = 7'h11 == _myNewVec_91_T_3[6:0] ? myVec_17 : _GEN_4794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4796 = 7'h12 == _myNewVec_91_T_3[6:0] ? myVec_18 : _GEN_4795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4797 = 7'h13 == _myNewVec_91_T_3[6:0] ? myVec_19 : _GEN_4796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4798 = 7'h14 == _myNewVec_91_T_3[6:0] ? myVec_20 : _GEN_4797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4799 = 7'h15 == _myNewVec_91_T_3[6:0] ? myVec_21 : _GEN_4798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4800 = 7'h16 == _myNewVec_91_T_3[6:0] ? myVec_22 : _GEN_4799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4801 = 7'h17 == _myNewVec_91_T_3[6:0] ? myVec_23 : _GEN_4800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4802 = 7'h18 == _myNewVec_91_T_3[6:0] ? myVec_24 : _GEN_4801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4803 = 7'h19 == _myNewVec_91_T_3[6:0] ? myVec_25 : _GEN_4802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4804 = 7'h1a == _myNewVec_91_T_3[6:0] ? myVec_26 : _GEN_4803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4805 = 7'h1b == _myNewVec_91_T_3[6:0] ? myVec_27 : _GEN_4804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4806 = 7'h1c == _myNewVec_91_T_3[6:0] ? myVec_28 : _GEN_4805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4807 = 7'h1d == _myNewVec_91_T_3[6:0] ? myVec_29 : _GEN_4806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4808 = 7'h1e == _myNewVec_91_T_3[6:0] ? myVec_30 : _GEN_4807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4809 = 7'h1f == _myNewVec_91_T_3[6:0] ? myVec_31 : _GEN_4808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4810 = 7'h20 == _myNewVec_91_T_3[6:0] ? myVec_32 : _GEN_4809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4811 = 7'h21 == _myNewVec_91_T_3[6:0] ? myVec_33 : _GEN_4810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4812 = 7'h22 == _myNewVec_91_T_3[6:0] ? myVec_34 : _GEN_4811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4813 = 7'h23 == _myNewVec_91_T_3[6:0] ? myVec_35 : _GEN_4812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4814 = 7'h24 == _myNewVec_91_T_3[6:0] ? myVec_36 : _GEN_4813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4815 = 7'h25 == _myNewVec_91_T_3[6:0] ? myVec_37 : _GEN_4814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4816 = 7'h26 == _myNewVec_91_T_3[6:0] ? myVec_38 : _GEN_4815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4817 = 7'h27 == _myNewVec_91_T_3[6:0] ? myVec_39 : _GEN_4816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4818 = 7'h28 == _myNewVec_91_T_3[6:0] ? myVec_40 : _GEN_4817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4819 = 7'h29 == _myNewVec_91_T_3[6:0] ? myVec_41 : _GEN_4818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4820 = 7'h2a == _myNewVec_91_T_3[6:0] ? myVec_42 : _GEN_4819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4821 = 7'h2b == _myNewVec_91_T_3[6:0] ? myVec_43 : _GEN_4820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4822 = 7'h2c == _myNewVec_91_T_3[6:0] ? myVec_44 : _GEN_4821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4823 = 7'h2d == _myNewVec_91_T_3[6:0] ? myVec_45 : _GEN_4822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4824 = 7'h2e == _myNewVec_91_T_3[6:0] ? myVec_46 : _GEN_4823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4825 = 7'h2f == _myNewVec_91_T_3[6:0] ? myVec_47 : _GEN_4824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4826 = 7'h30 == _myNewVec_91_T_3[6:0] ? myVec_48 : _GEN_4825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4827 = 7'h31 == _myNewVec_91_T_3[6:0] ? myVec_49 : _GEN_4826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4828 = 7'h32 == _myNewVec_91_T_3[6:0] ? myVec_50 : _GEN_4827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4829 = 7'h33 == _myNewVec_91_T_3[6:0] ? myVec_51 : _GEN_4828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4830 = 7'h34 == _myNewVec_91_T_3[6:0] ? myVec_52 : _GEN_4829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4831 = 7'h35 == _myNewVec_91_T_3[6:0] ? myVec_53 : _GEN_4830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4832 = 7'h36 == _myNewVec_91_T_3[6:0] ? myVec_54 : _GEN_4831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4833 = 7'h37 == _myNewVec_91_T_3[6:0] ? myVec_55 : _GEN_4832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4834 = 7'h38 == _myNewVec_91_T_3[6:0] ? myVec_56 : _GEN_4833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4835 = 7'h39 == _myNewVec_91_T_3[6:0] ? myVec_57 : _GEN_4834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4836 = 7'h3a == _myNewVec_91_T_3[6:0] ? myVec_58 : _GEN_4835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4837 = 7'h3b == _myNewVec_91_T_3[6:0] ? myVec_59 : _GEN_4836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4838 = 7'h3c == _myNewVec_91_T_3[6:0] ? myVec_60 : _GEN_4837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4839 = 7'h3d == _myNewVec_91_T_3[6:0] ? myVec_61 : _GEN_4838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4840 = 7'h3e == _myNewVec_91_T_3[6:0] ? myVec_62 : _GEN_4839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4841 = 7'h3f == _myNewVec_91_T_3[6:0] ? myVec_63 : _GEN_4840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4842 = 7'h40 == _myNewVec_91_T_3[6:0] ? myVec_64 : _GEN_4841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4843 = 7'h41 == _myNewVec_91_T_3[6:0] ? myVec_65 : _GEN_4842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4844 = 7'h42 == _myNewVec_91_T_3[6:0] ? myVec_66 : _GEN_4843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4845 = 7'h43 == _myNewVec_91_T_3[6:0] ? myVec_67 : _GEN_4844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4846 = 7'h44 == _myNewVec_91_T_3[6:0] ? myVec_68 : _GEN_4845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4847 = 7'h45 == _myNewVec_91_T_3[6:0] ? myVec_69 : _GEN_4846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4848 = 7'h46 == _myNewVec_91_T_3[6:0] ? myVec_70 : _GEN_4847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4849 = 7'h47 == _myNewVec_91_T_3[6:0] ? myVec_71 : _GEN_4848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4850 = 7'h48 == _myNewVec_91_T_3[6:0] ? myVec_72 : _GEN_4849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4851 = 7'h49 == _myNewVec_91_T_3[6:0] ? myVec_73 : _GEN_4850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4852 = 7'h4a == _myNewVec_91_T_3[6:0] ? myVec_74 : _GEN_4851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4853 = 7'h4b == _myNewVec_91_T_3[6:0] ? myVec_75 : _GEN_4852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4854 = 7'h4c == _myNewVec_91_T_3[6:0] ? myVec_76 : _GEN_4853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4855 = 7'h4d == _myNewVec_91_T_3[6:0] ? myVec_77 : _GEN_4854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4856 = 7'h4e == _myNewVec_91_T_3[6:0] ? myVec_78 : _GEN_4855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4857 = 7'h4f == _myNewVec_91_T_3[6:0] ? myVec_79 : _GEN_4856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4858 = 7'h50 == _myNewVec_91_T_3[6:0] ? myVec_80 : _GEN_4857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4859 = 7'h51 == _myNewVec_91_T_3[6:0] ? myVec_81 : _GEN_4858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4860 = 7'h52 == _myNewVec_91_T_3[6:0] ? myVec_82 : _GEN_4859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4861 = 7'h53 == _myNewVec_91_T_3[6:0] ? myVec_83 : _GEN_4860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4862 = 7'h54 == _myNewVec_91_T_3[6:0] ? myVec_84 : _GEN_4861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4863 = 7'h55 == _myNewVec_91_T_3[6:0] ? myVec_85 : _GEN_4862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4864 = 7'h56 == _myNewVec_91_T_3[6:0] ? myVec_86 : _GEN_4863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4865 = 7'h57 == _myNewVec_91_T_3[6:0] ? myVec_87 : _GEN_4864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4866 = 7'h58 == _myNewVec_91_T_3[6:0] ? myVec_88 : _GEN_4865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4867 = 7'h59 == _myNewVec_91_T_3[6:0] ? myVec_89 : _GEN_4866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4868 = 7'h5a == _myNewVec_91_T_3[6:0] ? myVec_90 : _GEN_4867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4869 = 7'h5b == _myNewVec_91_T_3[6:0] ? myVec_91 : _GEN_4868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4870 = 7'h5c == _myNewVec_91_T_3[6:0] ? myVec_92 : _GEN_4869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4871 = 7'h5d == _myNewVec_91_T_3[6:0] ? myVec_93 : _GEN_4870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4872 = 7'h5e == _myNewVec_91_T_3[6:0] ? myVec_94 : _GEN_4871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4873 = 7'h5f == _myNewVec_91_T_3[6:0] ? myVec_95 : _GEN_4872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4874 = 7'h60 == _myNewVec_91_T_3[6:0] ? myVec_96 : _GEN_4873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4875 = 7'h61 == _myNewVec_91_T_3[6:0] ? myVec_97 : _GEN_4874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4876 = 7'h62 == _myNewVec_91_T_3[6:0] ? myVec_98 : _GEN_4875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4877 = 7'h63 == _myNewVec_91_T_3[6:0] ? myVec_99 : _GEN_4876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4878 = 7'h64 == _myNewVec_91_T_3[6:0] ? myVec_100 : _GEN_4877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4879 = 7'h65 == _myNewVec_91_T_3[6:0] ? myVec_101 : _GEN_4878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4880 = 7'h66 == _myNewVec_91_T_3[6:0] ? myVec_102 : _GEN_4879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4881 = 7'h67 == _myNewVec_91_T_3[6:0] ? myVec_103 : _GEN_4880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4882 = 7'h68 == _myNewVec_91_T_3[6:0] ? myVec_104 : _GEN_4881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4883 = 7'h69 == _myNewVec_91_T_3[6:0] ? myVec_105 : _GEN_4882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4884 = 7'h6a == _myNewVec_91_T_3[6:0] ? myVec_106 : _GEN_4883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4885 = 7'h6b == _myNewVec_91_T_3[6:0] ? myVec_107 : _GEN_4884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4886 = 7'h6c == _myNewVec_91_T_3[6:0] ? myVec_108 : _GEN_4885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4887 = 7'h6d == _myNewVec_91_T_3[6:0] ? myVec_109 : _GEN_4886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4888 = 7'h6e == _myNewVec_91_T_3[6:0] ? myVec_110 : _GEN_4887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4889 = 7'h6f == _myNewVec_91_T_3[6:0] ? myVec_111 : _GEN_4888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4890 = 7'h70 == _myNewVec_91_T_3[6:0] ? myVec_112 : _GEN_4889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4891 = 7'h71 == _myNewVec_91_T_3[6:0] ? myVec_113 : _GEN_4890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4892 = 7'h72 == _myNewVec_91_T_3[6:0] ? myVec_114 : _GEN_4891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4893 = 7'h73 == _myNewVec_91_T_3[6:0] ? myVec_115 : _GEN_4892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4894 = 7'h74 == _myNewVec_91_T_3[6:0] ? myVec_116 : _GEN_4893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4895 = 7'h75 == _myNewVec_91_T_3[6:0] ? myVec_117 : _GEN_4894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4896 = 7'h76 == _myNewVec_91_T_3[6:0] ? myVec_118 : _GEN_4895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4897 = 7'h77 == _myNewVec_91_T_3[6:0] ? myVec_119 : _GEN_4896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4898 = 7'h78 == _myNewVec_91_T_3[6:0] ? myVec_120 : _GEN_4897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4899 = 7'h79 == _myNewVec_91_T_3[6:0] ? myVec_121 : _GEN_4898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4900 = 7'h7a == _myNewVec_91_T_3[6:0] ? myVec_122 : _GEN_4899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4901 = 7'h7b == _myNewVec_91_T_3[6:0] ? myVec_123 : _GEN_4900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4902 = 7'h7c == _myNewVec_91_T_3[6:0] ? myVec_124 : _GEN_4901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4903 = 7'h7d == _myNewVec_91_T_3[6:0] ? myVec_125 : _GEN_4902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4904 = 7'h7e == _myNewVec_91_T_3[6:0] ? myVec_126 : _GEN_4903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_91 = 7'h7f == _myNewVec_91_T_3[6:0] ? myVec_127 : _GEN_4904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_90_T_3 = _myNewVec_127_T_1 + 16'h25; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_4907 = 7'h1 == _myNewVec_90_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4908 = 7'h2 == _myNewVec_90_T_3[6:0] ? myVec_2 : _GEN_4907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4909 = 7'h3 == _myNewVec_90_T_3[6:0] ? myVec_3 : _GEN_4908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4910 = 7'h4 == _myNewVec_90_T_3[6:0] ? myVec_4 : _GEN_4909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4911 = 7'h5 == _myNewVec_90_T_3[6:0] ? myVec_5 : _GEN_4910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4912 = 7'h6 == _myNewVec_90_T_3[6:0] ? myVec_6 : _GEN_4911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4913 = 7'h7 == _myNewVec_90_T_3[6:0] ? myVec_7 : _GEN_4912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4914 = 7'h8 == _myNewVec_90_T_3[6:0] ? myVec_8 : _GEN_4913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4915 = 7'h9 == _myNewVec_90_T_3[6:0] ? myVec_9 : _GEN_4914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4916 = 7'ha == _myNewVec_90_T_3[6:0] ? myVec_10 : _GEN_4915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4917 = 7'hb == _myNewVec_90_T_3[6:0] ? myVec_11 : _GEN_4916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4918 = 7'hc == _myNewVec_90_T_3[6:0] ? myVec_12 : _GEN_4917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4919 = 7'hd == _myNewVec_90_T_3[6:0] ? myVec_13 : _GEN_4918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4920 = 7'he == _myNewVec_90_T_3[6:0] ? myVec_14 : _GEN_4919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4921 = 7'hf == _myNewVec_90_T_3[6:0] ? myVec_15 : _GEN_4920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4922 = 7'h10 == _myNewVec_90_T_3[6:0] ? myVec_16 : _GEN_4921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4923 = 7'h11 == _myNewVec_90_T_3[6:0] ? myVec_17 : _GEN_4922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4924 = 7'h12 == _myNewVec_90_T_3[6:0] ? myVec_18 : _GEN_4923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4925 = 7'h13 == _myNewVec_90_T_3[6:0] ? myVec_19 : _GEN_4924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4926 = 7'h14 == _myNewVec_90_T_3[6:0] ? myVec_20 : _GEN_4925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4927 = 7'h15 == _myNewVec_90_T_3[6:0] ? myVec_21 : _GEN_4926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4928 = 7'h16 == _myNewVec_90_T_3[6:0] ? myVec_22 : _GEN_4927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4929 = 7'h17 == _myNewVec_90_T_3[6:0] ? myVec_23 : _GEN_4928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4930 = 7'h18 == _myNewVec_90_T_3[6:0] ? myVec_24 : _GEN_4929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4931 = 7'h19 == _myNewVec_90_T_3[6:0] ? myVec_25 : _GEN_4930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4932 = 7'h1a == _myNewVec_90_T_3[6:0] ? myVec_26 : _GEN_4931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4933 = 7'h1b == _myNewVec_90_T_3[6:0] ? myVec_27 : _GEN_4932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4934 = 7'h1c == _myNewVec_90_T_3[6:0] ? myVec_28 : _GEN_4933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4935 = 7'h1d == _myNewVec_90_T_3[6:0] ? myVec_29 : _GEN_4934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4936 = 7'h1e == _myNewVec_90_T_3[6:0] ? myVec_30 : _GEN_4935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4937 = 7'h1f == _myNewVec_90_T_3[6:0] ? myVec_31 : _GEN_4936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4938 = 7'h20 == _myNewVec_90_T_3[6:0] ? myVec_32 : _GEN_4937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4939 = 7'h21 == _myNewVec_90_T_3[6:0] ? myVec_33 : _GEN_4938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4940 = 7'h22 == _myNewVec_90_T_3[6:0] ? myVec_34 : _GEN_4939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4941 = 7'h23 == _myNewVec_90_T_3[6:0] ? myVec_35 : _GEN_4940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4942 = 7'h24 == _myNewVec_90_T_3[6:0] ? myVec_36 : _GEN_4941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4943 = 7'h25 == _myNewVec_90_T_3[6:0] ? myVec_37 : _GEN_4942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4944 = 7'h26 == _myNewVec_90_T_3[6:0] ? myVec_38 : _GEN_4943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4945 = 7'h27 == _myNewVec_90_T_3[6:0] ? myVec_39 : _GEN_4944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4946 = 7'h28 == _myNewVec_90_T_3[6:0] ? myVec_40 : _GEN_4945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4947 = 7'h29 == _myNewVec_90_T_3[6:0] ? myVec_41 : _GEN_4946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4948 = 7'h2a == _myNewVec_90_T_3[6:0] ? myVec_42 : _GEN_4947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4949 = 7'h2b == _myNewVec_90_T_3[6:0] ? myVec_43 : _GEN_4948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4950 = 7'h2c == _myNewVec_90_T_3[6:0] ? myVec_44 : _GEN_4949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4951 = 7'h2d == _myNewVec_90_T_3[6:0] ? myVec_45 : _GEN_4950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4952 = 7'h2e == _myNewVec_90_T_3[6:0] ? myVec_46 : _GEN_4951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4953 = 7'h2f == _myNewVec_90_T_3[6:0] ? myVec_47 : _GEN_4952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4954 = 7'h30 == _myNewVec_90_T_3[6:0] ? myVec_48 : _GEN_4953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4955 = 7'h31 == _myNewVec_90_T_3[6:0] ? myVec_49 : _GEN_4954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4956 = 7'h32 == _myNewVec_90_T_3[6:0] ? myVec_50 : _GEN_4955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4957 = 7'h33 == _myNewVec_90_T_3[6:0] ? myVec_51 : _GEN_4956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4958 = 7'h34 == _myNewVec_90_T_3[6:0] ? myVec_52 : _GEN_4957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4959 = 7'h35 == _myNewVec_90_T_3[6:0] ? myVec_53 : _GEN_4958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4960 = 7'h36 == _myNewVec_90_T_3[6:0] ? myVec_54 : _GEN_4959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4961 = 7'h37 == _myNewVec_90_T_3[6:0] ? myVec_55 : _GEN_4960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4962 = 7'h38 == _myNewVec_90_T_3[6:0] ? myVec_56 : _GEN_4961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4963 = 7'h39 == _myNewVec_90_T_3[6:0] ? myVec_57 : _GEN_4962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4964 = 7'h3a == _myNewVec_90_T_3[6:0] ? myVec_58 : _GEN_4963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4965 = 7'h3b == _myNewVec_90_T_3[6:0] ? myVec_59 : _GEN_4964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4966 = 7'h3c == _myNewVec_90_T_3[6:0] ? myVec_60 : _GEN_4965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4967 = 7'h3d == _myNewVec_90_T_3[6:0] ? myVec_61 : _GEN_4966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4968 = 7'h3e == _myNewVec_90_T_3[6:0] ? myVec_62 : _GEN_4967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4969 = 7'h3f == _myNewVec_90_T_3[6:0] ? myVec_63 : _GEN_4968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4970 = 7'h40 == _myNewVec_90_T_3[6:0] ? myVec_64 : _GEN_4969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4971 = 7'h41 == _myNewVec_90_T_3[6:0] ? myVec_65 : _GEN_4970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4972 = 7'h42 == _myNewVec_90_T_3[6:0] ? myVec_66 : _GEN_4971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4973 = 7'h43 == _myNewVec_90_T_3[6:0] ? myVec_67 : _GEN_4972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4974 = 7'h44 == _myNewVec_90_T_3[6:0] ? myVec_68 : _GEN_4973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4975 = 7'h45 == _myNewVec_90_T_3[6:0] ? myVec_69 : _GEN_4974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4976 = 7'h46 == _myNewVec_90_T_3[6:0] ? myVec_70 : _GEN_4975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4977 = 7'h47 == _myNewVec_90_T_3[6:0] ? myVec_71 : _GEN_4976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4978 = 7'h48 == _myNewVec_90_T_3[6:0] ? myVec_72 : _GEN_4977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4979 = 7'h49 == _myNewVec_90_T_3[6:0] ? myVec_73 : _GEN_4978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4980 = 7'h4a == _myNewVec_90_T_3[6:0] ? myVec_74 : _GEN_4979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4981 = 7'h4b == _myNewVec_90_T_3[6:0] ? myVec_75 : _GEN_4980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4982 = 7'h4c == _myNewVec_90_T_3[6:0] ? myVec_76 : _GEN_4981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4983 = 7'h4d == _myNewVec_90_T_3[6:0] ? myVec_77 : _GEN_4982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4984 = 7'h4e == _myNewVec_90_T_3[6:0] ? myVec_78 : _GEN_4983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4985 = 7'h4f == _myNewVec_90_T_3[6:0] ? myVec_79 : _GEN_4984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4986 = 7'h50 == _myNewVec_90_T_3[6:0] ? myVec_80 : _GEN_4985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4987 = 7'h51 == _myNewVec_90_T_3[6:0] ? myVec_81 : _GEN_4986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4988 = 7'h52 == _myNewVec_90_T_3[6:0] ? myVec_82 : _GEN_4987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4989 = 7'h53 == _myNewVec_90_T_3[6:0] ? myVec_83 : _GEN_4988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4990 = 7'h54 == _myNewVec_90_T_3[6:0] ? myVec_84 : _GEN_4989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4991 = 7'h55 == _myNewVec_90_T_3[6:0] ? myVec_85 : _GEN_4990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4992 = 7'h56 == _myNewVec_90_T_3[6:0] ? myVec_86 : _GEN_4991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4993 = 7'h57 == _myNewVec_90_T_3[6:0] ? myVec_87 : _GEN_4992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4994 = 7'h58 == _myNewVec_90_T_3[6:0] ? myVec_88 : _GEN_4993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4995 = 7'h59 == _myNewVec_90_T_3[6:0] ? myVec_89 : _GEN_4994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4996 = 7'h5a == _myNewVec_90_T_3[6:0] ? myVec_90 : _GEN_4995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4997 = 7'h5b == _myNewVec_90_T_3[6:0] ? myVec_91 : _GEN_4996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4998 = 7'h5c == _myNewVec_90_T_3[6:0] ? myVec_92 : _GEN_4997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4999 = 7'h5d == _myNewVec_90_T_3[6:0] ? myVec_93 : _GEN_4998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5000 = 7'h5e == _myNewVec_90_T_3[6:0] ? myVec_94 : _GEN_4999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5001 = 7'h5f == _myNewVec_90_T_3[6:0] ? myVec_95 : _GEN_5000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5002 = 7'h60 == _myNewVec_90_T_3[6:0] ? myVec_96 : _GEN_5001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5003 = 7'h61 == _myNewVec_90_T_3[6:0] ? myVec_97 : _GEN_5002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5004 = 7'h62 == _myNewVec_90_T_3[6:0] ? myVec_98 : _GEN_5003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5005 = 7'h63 == _myNewVec_90_T_3[6:0] ? myVec_99 : _GEN_5004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5006 = 7'h64 == _myNewVec_90_T_3[6:0] ? myVec_100 : _GEN_5005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5007 = 7'h65 == _myNewVec_90_T_3[6:0] ? myVec_101 : _GEN_5006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5008 = 7'h66 == _myNewVec_90_T_3[6:0] ? myVec_102 : _GEN_5007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5009 = 7'h67 == _myNewVec_90_T_3[6:0] ? myVec_103 : _GEN_5008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5010 = 7'h68 == _myNewVec_90_T_3[6:0] ? myVec_104 : _GEN_5009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5011 = 7'h69 == _myNewVec_90_T_3[6:0] ? myVec_105 : _GEN_5010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5012 = 7'h6a == _myNewVec_90_T_3[6:0] ? myVec_106 : _GEN_5011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5013 = 7'h6b == _myNewVec_90_T_3[6:0] ? myVec_107 : _GEN_5012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5014 = 7'h6c == _myNewVec_90_T_3[6:0] ? myVec_108 : _GEN_5013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5015 = 7'h6d == _myNewVec_90_T_3[6:0] ? myVec_109 : _GEN_5014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5016 = 7'h6e == _myNewVec_90_T_3[6:0] ? myVec_110 : _GEN_5015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5017 = 7'h6f == _myNewVec_90_T_3[6:0] ? myVec_111 : _GEN_5016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5018 = 7'h70 == _myNewVec_90_T_3[6:0] ? myVec_112 : _GEN_5017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5019 = 7'h71 == _myNewVec_90_T_3[6:0] ? myVec_113 : _GEN_5018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5020 = 7'h72 == _myNewVec_90_T_3[6:0] ? myVec_114 : _GEN_5019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5021 = 7'h73 == _myNewVec_90_T_3[6:0] ? myVec_115 : _GEN_5020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5022 = 7'h74 == _myNewVec_90_T_3[6:0] ? myVec_116 : _GEN_5021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5023 = 7'h75 == _myNewVec_90_T_3[6:0] ? myVec_117 : _GEN_5022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5024 = 7'h76 == _myNewVec_90_T_3[6:0] ? myVec_118 : _GEN_5023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5025 = 7'h77 == _myNewVec_90_T_3[6:0] ? myVec_119 : _GEN_5024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5026 = 7'h78 == _myNewVec_90_T_3[6:0] ? myVec_120 : _GEN_5025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5027 = 7'h79 == _myNewVec_90_T_3[6:0] ? myVec_121 : _GEN_5026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5028 = 7'h7a == _myNewVec_90_T_3[6:0] ? myVec_122 : _GEN_5027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5029 = 7'h7b == _myNewVec_90_T_3[6:0] ? myVec_123 : _GEN_5028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5030 = 7'h7c == _myNewVec_90_T_3[6:0] ? myVec_124 : _GEN_5029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5031 = 7'h7d == _myNewVec_90_T_3[6:0] ? myVec_125 : _GEN_5030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5032 = 7'h7e == _myNewVec_90_T_3[6:0] ? myVec_126 : _GEN_5031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_90 = 7'h7f == _myNewVec_90_T_3[6:0] ? myVec_127 : _GEN_5032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_89_T_3 = _myNewVec_127_T_1 + 16'h26; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_5035 = 7'h1 == _myNewVec_89_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5036 = 7'h2 == _myNewVec_89_T_3[6:0] ? myVec_2 : _GEN_5035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5037 = 7'h3 == _myNewVec_89_T_3[6:0] ? myVec_3 : _GEN_5036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5038 = 7'h4 == _myNewVec_89_T_3[6:0] ? myVec_4 : _GEN_5037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5039 = 7'h5 == _myNewVec_89_T_3[6:0] ? myVec_5 : _GEN_5038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5040 = 7'h6 == _myNewVec_89_T_3[6:0] ? myVec_6 : _GEN_5039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5041 = 7'h7 == _myNewVec_89_T_3[6:0] ? myVec_7 : _GEN_5040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5042 = 7'h8 == _myNewVec_89_T_3[6:0] ? myVec_8 : _GEN_5041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5043 = 7'h9 == _myNewVec_89_T_3[6:0] ? myVec_9 : _GEN_5042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5044 = 7'ha == _myNewVec_89_T_3[6:0] ? myVec_10 : _GEN_5043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5045 = 7'hb == _myNewVec_89_T_3[6:0] ? myVec_11 : _GEN_5044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5046 = 7'hc == _myNewVec_89_T_3[6:0] ? myVec_12 : _GEN_5045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5047 = 7'hd == _myNewVec_89_T_3[6:0] ? myVec_13 : _GEN_5046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5048 = 7'he == _myNewVec_89_T_3[6:0] ? myVec_14 : _GEN_5047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5049 = 7'hf == _myNewVec_89_T_3[6:0] ? myVec_15 : _GEN_5048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5050 = 7'h10 == _myNewVec_89_T_3[6:0] ? myVec_16 : _GEN_5049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5051 = 7'h11 == _myNewVec_89_T_3[6:0] ? myVec_17 : _GEN_5050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5052 = 7'h12 == _myNewVec_89_T_3[6:0] ? myVec_18 : _GEN_5051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5053 = 7'h13 == _myNewVec_89_T_3[6:0] ? myVec_19 : _GEN_5052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5054 = 7'h14 == _myNewVec_89_T_3[6:0] ? myVec_20 : _GEN_5053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5055 = 7'h15 == _myNewVec_89_T_3[6:0] ? myVec_21 : _GEN_5054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5056 = 7'h16 == _myNewVec_89_T_3[6:0] ? myVec_22 : _GEN_5055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5057 = 7'h17 == _myNewVec_89_T_3[6:0] ? myVec_23 : _GEN_5056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5058 = 7'h18 == _myNewVec_89_T_3[6:0] ? myVec_24 : _GEN_5057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5059 = 7'h19 == _myNewVec_89_T_3[6:0] ? myVec_25 : _GEN_5058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5060 = 7'h1a == _myNewVec_89_T_3[6:0] ? myVec_26 : _GEN_5059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5061 = 7'h1b == _myNewVec_89_T_3[6:0] ? myVec_27 : _GEN_5060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5062 = 7'h1c == _myNewVec_89_T_3[6:0] ? myVec_28 : _GEN_5061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5063 = 7'h1d == _myNewVec_89_T_3[6:0] ? myVec_29 : _GEN_5062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5064 = 7'h1e == _myNewVec_89_T_3[6:0] ? myVec_30 : _GEN_5063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5065 = 7'h1f == _myNewVec_89_T_3[6:0] ? myVec_31 : _GEN_5064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5066 = 7'h20 == _myNewVec_89_T_3[6:0] ? myVec_32 : _GEN_5065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5067 = 7'h21 == _myNewVec_89_T_3[6:0] ? myVec_33 : _GEN_5066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5068 = 7'h22 == _myNewVec_89_T_3[6:0] ? myVec_34 : _GEN_5067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5069 = 7'h23 == _myNewVec_89_T_3[6:0] ? myVec_35 : _GEN_5068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5070 = 7'h24 == _myNewVec_89_T_3[6:0] ? myVec_36 : _GEN_5069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5071 = 7'h25 == _myNewVec_89_T_3[6:0] ? myVec_37 : _GEN_5070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5072 = 7'h26 == _myNewVec_89_T_3[6:0] ? myVec_38 : _GEN_5071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5073 = 7'h27 == _myNewVec_89_T_3[6:0] ? myVec_39 : _GEN_5072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5074 = 7'h28 == _myNewVec_89_T_3[6:0] ? myVec_40 : _GEN_5073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5075 = 7'h29 == _myNewVec_89_T_3[6:0] ? myVec_41 : _GEN_5074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5076 = 7'h2a == _myNewVec_89_T_3[6:0] ? myVec_42 : _GEN_5075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5077 = 7'h2b == _myNewVec_89_T_3[6:0] ? myVec_43 : _GEN_5076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5078 = 7'h2c == _myNewVec_89_T_3[6:0] ? myVec_44 : _GEN_5077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5079 = 7'h2d == _myNewVec_89_T_3[6:0] ? myVec_45 : _GEN_5078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5080 = 7'h2e == _myNewVec_89_T_3[6:0] ? myVec_46 : _GEN_5079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5081 = 7'h2f == _myNewVec_89_T_3[6:0] ? myVec_47 : _GEN_5080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5082 = 7'h30 == _myNewVec_89_T_3[6:0] ? myVec_48 : _GEN_5081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5083 = 7'h31 == _myNewVec_89_T_3[6:0] ? myVec_49 : _GEN_5082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5084 = 7'h32 == _myNewVec_89_T_3[6:0] ? myVec_50 : _GEN_5083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5085 = 7'h33 == _myNewVec_89_T_3[6:0] ? myVec_51 : _GEN_5084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5086 = 7'h34 == _myNewVec_89_T_3[6:0] ? myVec_52 : _GEN_5085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5087 = 7'h35 == _myNewVec_89_T_3[6:0] ? myVec_53 : _GEN_5086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5088 = 7'h36 == _myNewVec_89_T_3[6:0] ? myVec_54 : _GEN_5087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5089 = 7'h37 == _myNewVec_89_T_3[6:0] ? myVec_55 : _GEN_5088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5090 = 7'h38 == _myNewVec_89_T_3[6:0] ? myVec_56 : _GEN_5089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5091 = 7'h39 == _myNewVec_89_T_3[6:0] ? myVec_57 : _GEN_5090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5092 = 7'h3a == _myNewVec_89_T_3[6:0] ? myVec_58 : _GEN_5091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5093 = 7'h3b == _myNewVec_89_T_3[6:0] ? myVec_59 : _GEN_5092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5094 = 7'h3c == _myNewVec_89_T_3[6:0] ? myVec_60 : _GEN_5093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5095 = 7'h3d == _myNewVec_89_T_3[6:0] ? myVec_61 : _GEN_5094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5096 = 7'h3e == _myNewVec_89_T_3[6:0] ? myVec_62 : _GEN_5095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5097 = 7'h3f == _myNewVec_89_T_3[6:0] ? myVec_63 : _GEN_5096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5098 = 7'h40 == _myNewVec_89_T_3[6:0] ? myVec_64 : _GEN_5097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5099 = 7'h41 == _myNewVec_89_T_3[6:0] ? myVec_65 : _GEN_5098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5100 = 7'h42 == _myNewVec_89_T_3[6:0] ? myVec_66 : _GEN_5099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5101 = 7'h43 == _myNewVec_89_T_3[6:0] ? myVec_67 : _GEN_5100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5102 = 7'h44 == _myNewVec_89_T_3[6:0] ? myVec_68 : _GEN_5101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5103 = 7'h45 == _myNewVec_89_T_3[6:0] ? myVec_69 : _GEN_5102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5104 = 7'h46 == _myNewVec_89_T_3[6:0] ? myVec_70 : _GEN_5103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5105 = 7'h47 == _myNewVec_89_T_3[6:0] ? myVec_71 : _GEN_5104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5106 = 7'h48 == _myNewVec_89_T_3[6:0] ? myVec_72 : _GEN_5105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5107 = 7'h49 == _myNewVec_89_T_3[6:0] ? myVec_73 : _GEN_5106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5108 = 7'h4a == _myNewVec_89_T_3[6:0] ? myVec_74 : _GEN_5107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5109 = 7'h4b == _myNewVec_89_T_3[6:0] ? myVec_75 : _GEN_5108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5110 = 7'h4c == _myNewVec_89_T_3[6:0] ? myVec_76 : _GEN_5109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5111 = 7'h4d == _myNewVec_89_T_3[6:0] ? myVec_77 : _GEN_5110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5112 = 7'h4e == _myNewVec_89_T_3[6:0] ? myVec_78 : _GEN_5111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5113 = 7'h4f == _myNewVec_89_T_3[6:0] ? myVec_79 : _GEN_5112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5114 = 7'h50 == _myNewVec_89_T_3[6:0] ? myVec_80 : _GEN_5113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5115 = 7'h51 == _myNewVec_89_T_3[6:0] ? myVec_81 : _GEN_5114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5116 = 7'h52 == _myNewVec_89_T_3[6:0] ? myVec_82 : _GEN_5115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5117 = 7'h53 == _myNewVec_89_T_3[6:0] ? myVec_83 : _GEN_5116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5118 = 7'h54 == _myNewVec_89_T_3[6:0] ? myVec_84 : _GEN_5117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5119 = 7'h55 == _myNewVec_89_T_3[6:0] ? myVec_85 : _GEN_5118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5120 = 7'h56 == _myNewVec_89_T_3[6:0] ? myVec_86 : _GEN_5119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5121 = 7'h57 == _myNewVec_89_T_3[6:0] ? myVec_87 : _GEN_5120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5122 = 7'h58 == _myNewVec_89_T_3[6:0] ? myVec_88 : _GEN_5121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5123 = 7'h59 == _myNewVec_89_T_3[6:0] ? myVec_89 : _GEN_5122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5124 = 7'h5a == _myNewVec_89_T_3[6:0] ? myVec_90 : _GEN_5123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5125 = 7'h5b == _myNewVec_89_T_3[6:0] ? myVec_91 : _GEN_5124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5126 = 7'h5c == _myNewVec_89_T_3[6:0] ? myVec_92 : _GEN_5125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5127 = 7'h5d == _myNewVec_89_T_3[6:0] ? myVec_93 : _GEN_5126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5128 = 7'h5e == _myNewVec_89_T_3[6:0] ? myVec_94 : _GEN_5127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5129 = 7'h5f == _myNewVec_89_T_3[6:0] ? myVec_95 : _GEN_5128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5130 = 7'h60 == _myNewVec_89_T_3[6:0] ? myVec_96 : _GEN_5129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5131 = 7'h61 == _myNewVec_89_T_3[6:0] ? myVec_97 : _GEN_5130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5132 = 7'h62 == _myNewVec_89_T_3[6:0] ? myVec_98 : _GEN_5131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5133 = 7'h63 == _myNewVec_89_T_3[6:0] ? myVec_99 : _GEN_5132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5134 = 7'h64 == _myNewVec_89_T_3[6:0] ? myVec_100 : _GEN_5133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5135 = 7'h65 == _myNewVec_89_T_3[6:0] ? myVec_101 : _GEN_5134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5136 = 7'h66 == _myNewVec_89_T_3[6:0] ? myVec_102 : _GEN_5135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5137 = 7'h67 == _myNewVec_89_T_3[6:0] ? myVec_103 : _GEN_5136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5138 = 7'h68 == _myNewVec_89_T_3[6:0] ? myVec_104 : _GEN_5137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5139 = 7'h69 == _myNewVec_89_T_3[6:0] ? myVec_105 : _GEN_5138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5140 = 7'h6a == _myNewVec_89_T_3[6:0] ? myVec_106 : _GEN_5139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5141 = 7'h6b == _myNewVec_89_T_3[6:0] ? myVec_107 : _GEN_5140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5142 = 7'h6c == _myNewVec_89_T_3[6:0] ? myVec_108 : _GEN_5141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5143 = 7'h6d == _myNewVec_89_T_3[6:0] ? myVec_109 : _GEN_5142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5144 = 7'h6e == _myNewVec_89_T_3[6:0] ? myVec_110 : _GEN_5143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5145 = 7'h6f == _myNewVec_89_T_3[6:0] ? myVec_111 : _GEN_5144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5146 = 7'h70 == _myNewVec_89_T_3[6:0] ? myVec_112 : _GEN_5145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5147 = 7'h71 == _myNewVec_89_T_3[6:0] ? myVec_113 : _GEN_5146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5148 = 7'h72 == _myNewVec_89_T_3[6:0] ? myVec_114 : _GEN_5147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5149 = 7'h73 == _myNewVec_89_T_3[6:0] ? myVec_115 : _GEN_5148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5150 = 7'h74 == _myNewVec_89_T_3[6:0] ? myVec_116 : _GEN_5149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5151 = 7'h75 == _myNewVec_89_T_3[6:0] ? myVec_117 : _GEN_5150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5152 = 7'h76 == _myNewVec_89_T_3[6:0] ? myVec_118 : _GEN_5151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5153 = 7'h77 == _myNewVec_89_T_3[6:0] ? myVec_119 : _GEN_5152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5154 = 7'h78 == _myNewVec_89_T_3[6:0] ? myVec_120 : _GEN_5153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5155 = 7'h79 == _myNewVec_89_T_3[6:0] ? myVec_121 : _GEN_5154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5156 = 7'h7a == _myNewVec_89_T_3[6:0] ? myVec_122 : _GEN_5155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5157 = 7'h7b == _myNewVec_89_T_3[6:0] ? myVec_123 : _GEN_5156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5158 = 7'h7c == _myNewVec_89_T_3[6:0] ? myVec_124 : _GEN_5157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5159 = 7'h7d == _myNewVec_89_T_3[6:0] ? myVec_125 : _GEN_5158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5160 = 7'h7e == _myNewVec_89_T_3[6:0] ? myVec_126 : _GEN_5159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_89 = 7'h7f == _myNewVec_89_T_3[6:0] ? myVec_127 : _GEN_5160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_88_T_3 = _myNewVec_127_T_1 + 16'h27; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_5163 = 7'h1 == _myNewVec_88_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5164 = 7'h2 == _myNewVec_88_T_3[6:0] ? myVec_2 : _GEN_5163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5165 = 7'h3 == _myNewVec_88_T_3[6:0] ? myVec_3 : _GEN_5164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5166 = 7'h4 == _myNewVec_88_T_3[6:0] ? myVec_4 : _GEN_5165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5167 = 7'h5 == _myNewVec_88_T_3[6:0] ? myVec_5 : _GEN_5166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5168 = 7'h6 == _myNewVec_88_T_3[6:0] ? myVec_6 : _GEN_5167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5169 = 7'h7 == _myNewVec_88_T_3[6:0] ? myVec_7 : _GEN_5168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5170 = 7'h8 == _myNewVec_88_T_3[6:0] ? myVec_8 : _GEN_5169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5171 = 7'h9 == _myNewVec_88_T_3[6:0] ? myVec_9 : _GEN_5170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5172 = 7'ha == _myNewVec_88_T_3[6:0] ? myVec_10 : _GEN_5171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5173 = 7'hb == _myNewVec_88_T_3[6:0] ? myVec_11 : _GEN_5172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5174 = 7'hc == _myNewVec_88_T_3[6:0] ? myVec_12 : _GEN_5173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5175 = 7'hd == _myNewVec_88_T_3[6:0] ? myVec_13 : _GEN_5174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5176 = 7'he == _myNewVec_88_T_3[6:0] ? myVec_14 : _GEN_5175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5177 = 7'hf == _myNewVec_88_T_3[6:0] ? myVec_15 : _GEN_5176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5178 = 7'h10 == _myNewVec_88_T_3[6:0] ? myVec_16 : _GEN_5177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5179 = 7'h11 == _myNewVec_88_T_3[6:0] ? myVec_17 : _GEN_5178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5180 = 7'h12 == _myNewVec_88_T_3[6:0] ? myVec_18 : _GEN_5179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5181 = 7'h13 == _myNewVec_88_T_3[6:0] ? myVec_19 : _GEN_5180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5182 = 7'h14 == _myNewVec_88_T_3[6:0] ? myVec_20 : _GEN_5181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5183 = 7'h15 == _myNewVec_88_T_3[6:0] ? myVec_21 : _GEN_5182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5184 = 7'h16 == _myNewVec_88_T_3[6:0] ? myVec_22 : _GEN_5183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5185 = 7'h17 == _myNewVec_88_T_3[6:0] ? myVec_23 : _GEN_5184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5186 = 7'h18 == _myNewVec_88_T_3[6:0] ? myVec_24 : _GEN_5185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5187 = 7'h19 == _myNewVec_88_T_3[6:0] ? myVec_25 : _GEN_5186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5188 = 7'h1a == _myNewVec_88_T_3[6:0] ? myVec_26 : _GEN_5187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5189 = 7'h1b == _myNewVec_88_T_3[6:0] ? myVec_27 : _GEN_5188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5190 = 7'h1c == _myNewVec_88_T_3[6:0] ? myVec_28 : _GEN_5189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5191 = 7'h1d == _myNewVec_88_T_3[6:0] ? myVec_29 : _GEN_5190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5192 = 7'h1e == _myNewVec_88_T_3[6:0] ? myVec_30 : _GEN_5191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5193 = 7'h1f == _myNewVec_88_T_3[6:0] ? myVec_31 : _GEN_5192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5194 = 7'h20 == _myNewVec_88_T_3[6:0] ? myVec_32 : _GEN_5193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5195 = 7'h21 == _myNewVec_88_T_3[6:0] ? myVec_33 : _GEN_5194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5196 = 7'h22 == _myNewVec_88_T_3[6:0] ? myVec_34 : _GEN_5195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5197 = 7'h23 == _myNewVec_88_T_3[6:0] ? myVec_35 : _GEN_5196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5198 = 7'h24 == _myNewVec_88_T_3[6:0] ? myVec_36 : _GEN_5197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5199 = 7'h25 == _myNewVec_88_T_3[6:0] ? myVec_37 : _GEN_5198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5200 = 7'h26 == _myNewVec_88_T_3[6:0] ? myVec_38 : _GEN_5199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5201 = 7'h27 == _myNewVec_88_T_3[6:0] ? myVec_39 : _GEN_5200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5202 = 7'h28 == _myNewVec_88_T_3[6:0] ? myVec_40 : _GEN_5201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5203 = 7'h29 == _myNewVec_88_T_3[6:0] ? myVec_41 : _GEN_5202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5204 = 7'h2a == _myNewVec_88_T_3[6:0] ? myVec_42 : _GEN_5203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5205 = 7'h2b == _myNewVec_88_T_3[6:0] ? myVec_43 : _GEN_5204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5206 = 7'h2c == _myNewVec_88_T_3[6:0] ? myVec_44 : _GEN_5205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5207 = 7'h2d == _myNewVec_88_T_3[6:0] ? myVec_45 : _GEN_5206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5208 = 7'h2e == _myNewVec_88_T_3[6:0] ? myVec_46 : _GEN_5207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5209 = 7'h2f == _myNewVec_88_T_3[6:0] ? myVec_47 : _GEN_5208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5210 = 7'h30 == _myNewVec_88_T_3[6:0] ? myVec_48 : _GEN_5209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5211 = 7'h31 == _myNewVec_88_T_3[6:0] ? myVec_49 : _GEN_5210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5212 = 7'h32 == _myNewVec_88_T_3[6:0] ? myVec_50 : _GEN_5211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5213 = 7'h33 == _myNewVec_88_T_3[6:0] ? myVec_51 : _GEN_5212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5214 = 7'h34 == _myNewVec_88_T_3[6:0] ? myVec_52 : _GEN_5213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5215 = 7'h35 == _myNewVec_88_T_3[6:0] ? myVec_53 : _GEN_5214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5216 = 7'h36 == _myNewVec_88_T_3[6:0] ? myVec_54 : _GEN_5215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5217 = 7'h37 == _myNewVec_88_T_3[6:0] ? myVec_55 : _GEN_5216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5218 = 7'h38 == _myNewVec_88_T_3[6:0] ? myVec_56 : _GEN_5217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5219 = 7'h39 == _myNewVec_88_T_3[6:0] ? myVec_57 : _GEN_5218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5220 = 7'h3a == _myNewVec_88_T_3[6:0] ? myVec_58 : _GEN_5219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5221 = 7'h3b == _myNewVec_88_T_3[6:0] ? myVec_59 : _GEN_5220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5222 = 7'h3c == _myNewVec_88_T_3[6:0] ? myVec_60 : _GEN_5221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5223 = 7'h3d == _myNewVec_88_T_3[6:0] ? myVec_61 : _GEN_5222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5224 = 7'h3e == _myNewVec_88_T_3[6:0] ? myVec_62 : _GEN_5223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5225 = 7'h3f == _myNewVec_88_T_3[6:0] ? myVec_63 : _GEN_5224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5226 = 7'h40 == _myNewVec_88_T_3[6:0] ? myVec_64 : _GEN_5225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5227 = 7'h41 == _myNewVec_88_T_3[6:0] ? myVec_65 : _GEN_5226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5228 = 7'h42 == _myNewVec_88_T_3[6:0] ? myVec_66 : _GEN_5227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5229 = 7'h43 == _myNewVec_88_T_3[6:0] ? myVec_67 : _GEN_5228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5230 = 7'h44 == _myNewVec_88_T_3[6:0] ? myVec_68 : _GEN_5229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5231 = 7'h45 == _myNewVec_88_T_3[6:0] ? myVec_69 : _GEN_5230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5232 = 7'h46 == _myNewVec_88_T_3[6:0] ? myVec_70 : _GEN_5231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5233 = 7'h47 == _myNewVec_88_T_3[6:0] ? myVec_71 : _GEN_5232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5234 = 7'h48 == _myNewVec_88_T_3[6:0] ? myVec_72 : _GEN_5233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5235 = 7'h49 == _myNewVec_88_T_3[6:0] ? myVec_73 : _GEN_5234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5236 = 7'h4a == _myNewVec_88_T_3[6:0] ? myVec_74 : _GEN_5235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5237 = 7'h4b == _myNewVec_88_T_3[6:0] ? myVec_75 : _GEN_5236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5238 = 7'h4c == _myNewVec_88_T_3[6:0] ? myVec_76 : _GEN_5237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5239 = 7'h4d == _myNewVec_88_T_3[6:0] ? myVec_77 : _GEN_5238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5240 = 7'h4e == _myNewVec_88_T_3[6:0] ? myVec_78 : _GEN_5239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5241 = 7'h4f == _myNewVec_88_T_3[6:0] ? myVec_79 : _GEN_5240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5242 = 7'h50 == _myNewVec_88_T_3[6:0] ? myVec_80 : _GEN_5241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5243 = 7'h51 == _myNewVec_88_T_3[6:0] ? myVec_81 : _GEN_5242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5244 = 7'h52 == _myNewVec_88_T_3[6:0] ? myVec_82 : _GEN_5243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5245 = 7'h53 == _myNewVec_88_T_3[6:0] ? myVec_83 : _GEN_5244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5246 = 7'h54 == _myNewVec_88_T_3[6:0] ? myVec_84 : _GEN_5245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5247 = 7'h55 == _myNewVec_88_T_3[6:0] ? myVec_85 : _GEN_5246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5248 = 7'h56 == _myNewVec_88_T_3[6:0] ? myVec_86 : _GEN_5247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5249 = 7'h57 == _myNewVec_88_T_3[6:0] ? myVec_87 : _GEN_5248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5250 = 7'h58 == _myNewVec_88_T_3[6:0] ? myVec_88 : _GEN_5249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5251 = 7'h59 == _myNewVec_88_T_3[6:0] ? myVec_89 : _GEN_5250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5252 = 7'h5a == _myNewVec_88_T_3[6:0] ? myVec_90 : _GEN_5251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5253 = 7'h5b == _myNewVec_88_T_3[6:0] ? myVec_91 : _GEN_5252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5254 = 7'h5c == _myNewVec_88_T_3[6:0] ? myVec_92 : _GEN_5253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5255 = 7'h5d == _myNewVec_88_T_3[6:0] ? myVec_93 : _GEN_5254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5256 = 7'h5e == _myNewVec_88_T_3[6:0] ? myVec_94 : _GEN_5255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5257 = 7'h5f == _myNewVec_88_T_3[6:0] ? myVec_95 : _GEN_5256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5258 = 7'h60 == _myNewVec_88_T_3[6:0] ? myVec_96 : _GEN_5257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5259 = 7'h61 == _myNewVec_88_T_3[6:0] ? myVec_97 : _GEN_5258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5260 = 7'h62 == _myNewVec_88_T_3[6:0] ? myVec_98 : _GEN_5259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5261 = 7'h63 == _myNewVec_88_T_3[6:0] ? myVec_99 : _GEN_5260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5262 = 7'h64 == _myNewVec_88_T_3[6:0] ? myVec_100 : _GEN_5261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5263 = 7'h65 == _myNewVec_88_T_3[6:0] ? myVec_101 : _GEN_5262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5264 = 7'h66 == _myNewVec_88_T_3[6:0] ? myVec_102 : _GEN_5263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5265 = 7'h67 == _myNewVec_88_T_3[6:0] ? myVec_103 : _GEN_5264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5266 = 7'h68 == _myNewVec_88_T_3[6:0] ? myVec_104 : _GEN_5265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5267 = 7'h69 == _myNewVec_88_T_3[6:0] ? myVec_105 : _GEN_5266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5268 = 7'h6a == _myNewVec_88_T_3[6:0] ? myVec_106 : _GEN_5267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5269 = 7'h6b == _myNewVec_88_T_3[6:0] ? myVec_107 : _GEN_5268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5270 = 7'h6c == _myNewVec_88_T_3[6:0] ? myVec_108 : _GEN_5269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5271 = 7'h6d == _myNewVec_88_T_3[6:0] ? myVec_109 : _GEN_5270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5272 = 7'h6e == _myNewVec_88_T_3[6:0] ? myVec_110 : _GEN_5271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5273 = 7'h6f == _myNewVec_88_T_3[6:0] ? myVec_111 : _GEN_5272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5274 = 7'h70 == _myNewVec_88_T_3[6:0] ? myVec_112 : _GEN_5273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5275 = 7'h71 == _myNewVec_88_T_3[6:0] ? myVec_113 : _GEN_5274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5276 = 7'h72 == _myNewVec_88_T_3[6:0] ? myVec_114 : _GEN_5275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5277 = 7'h73 == _myNewVec_88_T_3[6:0] ? myVec_115 : _GEN_5276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5278 = 7'h74 == _myNewVec_88_T_3[6:0] ? myVec_116 : _GEN_5277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5279 = 7'h75 == _myNewVec_88_T_3[6:0] ? myVec_117 : _GEN_5278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5280 = 7'h76 == _myNewVec_88_T_3[6:0] ? myVec_118 : _GEN_5279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5281 = 7'h77 == _myNewVec_88_T_3[6:0] ? myVec_119 : _GEN_5280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5282 = 7'h78 == _myNewVec_88_T_3[6:0] ? myVec_120 : _GEN_5281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5283 = 7'h79 == _myNewVec_88_T_3[6:0] ? myVec_121 : _GEN_5282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5284 = 7'h7a == _myNewVec_88_T_3[6:0] ? myVec_122 : _GEN_5283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5285 = 7'h7b == _myNewVec_88_T_3[6:0] ? myVec_123 : _GEN_5284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5286 = 7'h7c == _myNewVec_88_T_3[6:0] ? myVec_124 : _GEN_5285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5287 = 7'h7d == _myNewVec_88_T_3[6:0] ? myVec_125 : _GEN_5286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5288 = 7'h7e == _myNewVec_88_T_3[6:0] ? myVec_126 : _GEN_5287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_88 = 7'h7f == _myNewVec_88_T_3[6:0] ? myVec_127 : _GEN_5288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_87_T_3 = _myNewVec_127_T_1 + 16'h28; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_5291 = 7'h1 == _myNewVec_87_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5292 = 7'h2 == _myNewVec_87_T_3[6:0] ? myVec_2 : _GEN_5291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5293 = 7'h3 == _myNewVec_87_T_3[6:0] ? myVec_3 : _GEN_5292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5294 = 7'h4 == _myNewVec_87_T_3[6:0] ? myVec_4 : _GEN_5293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5295 = 7'h5 == _myNewVec_87_T_3[6:0] ? myVec_5 : _GEN_5294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5296 = 7'h6 == _myNewVec_87_T_3[6:0] ? myVec_6 : _GEN_5295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5297 = 7'h7 == _myNewVec_87_T_3[6:0] ? myVec_7 : _GEN_5296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5298 = 7'h8 == _myNewVec_87_T_3[6:0] ? myVec_8 : _GEN_5297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5299 = 7'h9 == _myNewVec_87_T_3[6:0] ? myVec_9 : _GEN_5298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5300 = 7'ha == _myNewVec_87_T_3[6:0] ? myVec_10 : _GEN_5299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5301 = 7'hb == _myNewVec_87_T_3[6:0] ? myVec_11 : _GEN_5300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5302 = 7'hc == _myNewVec_87_T_3[6:0] ? myVec_12 : _GEN_5301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5303 = 7'hd == _myNewVec_87_T_3[6:0] ? myVec_13 : _GEN_5302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5304 = 7'he == _myNewVec_87_T_3[6:0] ? myVec_14 : _GEN_5303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5305 = 7'hf == _myNewVec_87_T_3[6:0] ? myVec_15 : _GEN_5304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5306 = 7'h10 == _myNewVec_87_T_3[6:0] ? myVec_16 : _GEN_5305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5307 = 7'h11 == _myNewVec_87_T_3[6:0] ? myVec_17 : _GEN_5306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5308 = 7'h12 == _myNewVec_87_T_3[6:0] ? myVec_18 : _GEN_5307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5309 = 7'h13 == _myNewVec_87_T_3[6:0] ? myVec_19 : _GEN_5308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5310 = 7'h14 == _myNewVec_87_T_3[6:0] ? myVec_20 : _GEN_5309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5311 = 7'h15 == _myNewVec_87_T_3[6:0] ? myVec_21 : _GEN_5310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5312 = 7'h16 == _myNewVec_87_T_3[6:0] ? myVec_22 : _GEN_5311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5313 = 7'h17 == _myNewVec_87_T_3[6:0] ? myVec_23 : _GEN_5312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5314 = 7'h18 == _myNewVec_87_T_3[6:0] ? myVec_24 : _GEN_5313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5315 = 7'h19 == _myNewVec_87_T_3[6:0] ? myVec_25 : _GEN_5314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5316 = 7'h1a == _myNewVec_87_T_3[6:0] ? myVec_26 : _GEN_5315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5317 = 7'h1b == _myNewVec_87_T_3[6:0] ? myVec_27 : _GEN_5316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5318 = 7'h1c == _myNewVec_87_T_3[6:0] ? myVec_28 : _GEN_5317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5319 = 7'h1d == _myNewVec_87_T_3[6:0] ? myVec_29 : _GEN_5318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5320 = 7'h1e == _myNewVec_87_T_3[6:0] ? myVec_30 : _GEN_5319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5321 = 7'h1f == _myNewVec_87_T_3[6:0] ? myVec_31 : _GEN_5320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5322 = 7'h20 == _myNewVec_87_T_3[6:0] ? myVec_32 : _GEN_5321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5323 = 7'h21 == _myNewVec_87_T_3[6:0] ? myVec_33 : _GEN_5322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5324 = 7'h22 == _myNewVec_87_T_3[6:0] ? myVec_34 : _GEN_5323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5325 = 7'h23 == _myNewVec_87_T_3[6:0] ? myVec_35 : _GEN_5324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5326 = 7'h24 == _myNewVec_87_T_3[6:0] ? myVec_36 : _GEN_5325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5327 = 7'h25 == _myNewVec_87_T_3[6:0] ? myVec_37 : _GEN_5326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5328 = 7'h26 == _myNewVec_87_T_3[6:0] ? myVec_38 : _GEN_5327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5329 = 7'h27 == _myNewVec_87_T_3[6:0] ? myVec_39 : _GEN_5328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5330 = 7'h28 == _myNewVec_87_T_3[6:0] ? myVec_40 : _GEN_5329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5331 = 7'h29 == _myNewVec_87_T_3[6:0] ? myVec_41 : _GEN_5330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5332 = 7'h2a == _myNewVec_87_T_3[6:0] ? myVec_42 : _GEN_5331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5333 = 7'h2b == _myNewVec_87_T_3[6:0] ? myVec_43 : _GEN_5332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5334 = 7'h2c == _myNewVec_87_T_3[6:0] ? myVec_44 : _GEN_5333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5335 = 7'h2d == _myNewVec_87_T_3[6:0] ? myVec_45 : _GEN_5334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5336 = 7'h2e == _myNewVec_87_T_3[6:0] ? myVec_46 : _GEN_5335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5337 = 7'h2f == _myNewVec_87_T_3[6:0] ? myVec_47 : _GEN_5336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5338 = 7'h30 == _myNewVec_87_T_3[6:0] ? myVec_48 : _GEN_5337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5339 = 7'h31 == _myNewVec_87_T_3[6:0] ? myVec_49 : _GEN_5338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5340 = 7'h32 == _myNewVec_87_T_3[6:0] ? myVec_50 : _GEN_5339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5341 = 7'h33 == _myNewVec_87_T_3[6:0] ? myVec_51 : _GEN_5340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5342 = 7'h34 == _myNewVec_87_T_3[6:0] ? myVec_52 : _GEN_5341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5343 = 7'h35 == _myNewVec_87_T_3[6:0] ? myVec_53 : _GEN_5342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5344 = 7'h36 == _myNewVec_87_T_3[6:0] ? myVec_54 : _GEN_5343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5345 = 7'h37 == _myNewVec_87_T_3[6:0] ? myVec_55 : _GEN_5344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5346 = 7'h38 == _myNewVec_87_T_3[6:0] ? myVec_56 : _GEN_5345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5347 = 7'h39 == _myNewVec_87_T_3[6:0] ? myVec_57 : _GEN_5346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5348 = 7'h3a == _myNewVec_87_T_3[6:0] ? myVec_58 : _GEN_5347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5349 = 7'h3b == _myNewVec_87_T_3[6:0] ? myVec_59 : _GEN_5348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5350 = 7'h3c == _myNewVec_87_T_3[6:0] ? myVec_60 : _GEN_5349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5351 = 7'h3d == _myNewVec_87_T_3[6:0] ? myVec_61 : _GEN_5350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5352 = 7'h3e == _myNewVec_87_T_3[6:0] ? myVec_62 : _GEN_5351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5353 = 7'h3f == _myNewVec_87_T_3[6:0] ? myVec_63 : _GEN_5352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5354 = 7'h40 == _myNewVec_87_T_3[6:0] ? myVec_64 : _GEN_5353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5355 = 7'h41 == _myNewVec_87_T_3[6:0] ? myVec_65 : _GEN_5354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5356 = 7'h42 == _myNewVec_87_T_3[6:0] ? myVec_66 : _GEN_5355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5357 = 7'h43 == _myNewVec_87_T_3[6:0] ? myVec_67 : _GEN_5356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5358 = 7'h44 == _myNewVec_87_T_3[6:0] ? myVec_68 : _GEN_5357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5359 = 7'h45 == _myNewVec_87_T_3[6:0] ? myVec_69 : _GEN_5358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5360 = 7'h46 == _myNewVec_87_T_3[6:0] ? myVec_70 : _GEN_5359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5361 = 7'h47 == _myNewVec_87_T_3[6:0] ? myVec_71 : _GEN_5360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5362 = 7'h48 == _myNewVec_87_T_3[6:0] ? myVec_72 : _GEN_5361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5363 = 7'h49 == _myNewVec_87_T_3[6:0] ? myVec_73 : _GEN_5362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5364 = 7'h4a == _myNewVec_87_T_3[6:0] ? myVec_74 : _GEN_5363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5365 = 7'h4b == _myNewVec_87_T_3[6:0] ? myVec_75 : _GEN_5364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5366 = 7'h4c == _myNewVec_87_T_3[6:0] ? myVec_76 : _GEN_5365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5367 = 7'h4d == _myNewVec_87_T_3[6:0] ? myVec_77 : _GEN_5366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5368 = 7'h4e == _myNewVec_87_T_3[6:0] ? myVec_78 : _GEN_5367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5369 = 7'h4f == _myNewVec_87_T_3[6:0] ? myVec_79 : _GEN_5368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5370 = 7'h50 == _myNewVec_87_T_3[6:0] ? myVec_80 : _GEN_5369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5371 = 7'h51 == _myNewVec_87_T_3[6:0] ? myVec_81 : _GEN_5370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5372 = 7'h52 == _myNewVec_87_T_3[6:0] ? myVec_82 : _GEN_5371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5373 = 7'h53 == _myNewVec_87_T_3[6:0] ? myVec_83 : _GEN_5372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5374 = 7'h54 == _myNewVec_87_T_3[6:0] ? myVec_84 : _GEN_5373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5375 = 7'h55 == _myNewVec_87_T_3[6:0] ? myVec_85 : _GEN_5374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5376 = 7'h56 == _myNewVec_87_T_3[6:0] ? myVec_86 : _GEN_5375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5377 = 7'h57 == _myNewVec_87_T_3[6:0] ? myVec_87 : _GEN_5376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5378 = 7'h58 == _myNewVec_87_T_3[6:0] ? myVec_88 : _GEN_5377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5379 = 7'h59 == _myNewVec_87_T_3[6:0] ? myVec_89 : _GEN_5378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5380 = 7'h5a == _myNewVec_87_T_3[6:0] ? myVec_90 : _GEN_5379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5381 = 7'h5b == _myNewVec_87_T_3[6:0] ? myVec_91 : _GEN_5380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5382 = 7'h5c == _myNewVec_87_T_3[6:0] ? myVec_92 : _GEN_5381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5383 = 7'h5d == _myNewVec_87_T_3[6:0] ? myVec_93 : _GEN_5382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5384 = 7'h5e == _myNewVec_87_T_3[6:0] ? myVec_94 : _GEN_5383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5385 = 7'h5f == _myNewVec_87_T_3[6:0] ? myVec_95 : _GEN_5384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5386 = 7'h60 == _myNewVec_87_T_3[6:0] ? myVec_96 : _GEN_5385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5387 = 7'h61 == _myNewVec_87_T_3[6:0] ? myVec_97 : _GEN_5386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5388 = 7'h62 == _myNewVec_87_T_3[6:0] ? myVec_98 : _GEN_5387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5389 = 7'h63 == _myNewVec_87_T_3[6:0] ? myVec_99 : _GEN_5388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5390 = 7'h64 == _myNewVec_87_T_3[6:0] ? myVec_100 : _GEN_5389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5391 = 7'h65 == _myNewVec_87_T_3[6:0] ? myVec_101 : _GEN_5390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5392 = 7'h66 == _myNewVec_87_T_3[6:0] ? myVec_102 : _GEN_5391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5393 = 7'h67 == _myNewVec_87_T_3[6:0] ? myVec_103 : _GEN_5392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5394 = 7'h68 == _myNewVec_87_T_3[6:0] ? myVec_104 : _GEN_5393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5395 = 7'h69 == _myNewVec_87_T_3[6:0] ? myVec_105 : _GEN_5394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5396 = 7'h6a == _myNewVec_87_T_3[6:0] ? myVec_106 : _GEN_5395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5397 = 7'h6b == _myNewVec_87_T_3[6:0] ? myVec_107 : _GEN_5396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5398 = 7'h6c == _myNewVec_87_T_3[6:0] ? myVec_108 : _GEN_5397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5399 = 7'h6d == _myNewVec_87_T_3[6:0] ? myVec_109 : _GEN_5398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5400 = 7'h6e == _myNewVec_87_T_3[6:0] ? myVec_110 : _GEN_5399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5401 = 7'h6f == _myNewVec_87_T_3[6:0] ? myVec_111 : _GEN_5400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5402 = 7'h70 == _myNewVec_87_T_3[6:0] ? myVec_112 : _GEN_5401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5403 = 7'h71 == _myNewVec_87_T_3[6:0] ? myVec_113 : _GEN_5402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5404 = 7'h72 == _myNewVec_87_T_3[6:0] ? myVec_114 : _GEN_5403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5405 = 7'h73 == _myNewVec_87_T_3[6:0] ? myVec_115 : _GEN_5404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5406 = 7'h74 == _myNewVec_87_T_3[6:0] ? myVec_116 : _GEN_5405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5407 = 7'h75 == _myNewVec_87_T_3[6:0] ? myVec_117 : _GEN_5406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5408 = 7'h76 == _myNewVec_87_T_3[6:0] ? myVec_118 : _GEN_5407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5409 = 7'h77 == _myNewVec_87_T_3[6:0] ? myVec_119 : _GEN_5408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5410 = 7'h78 == _myNewVec_87_T_3[6:0] ? myVec_120 : _GEN_5409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5411 = 7'h79 == _myNewVec_87_T_3[6:0] ? myVec_121 : _GEN_5410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5412 = 7'h7a == _myNewVec_87_T_3[6:0] ? myVec_122 : _GEN_5411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5413 = 7'h7b == _myNewVec_87_T_3[6:0] ? myVec_123 : _GEN_5412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5414 = 7'h7c == _myNewVec_87_T_3[6:0] ? myVec_124 : _GEN_5413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5415 = 7'h7d == _myNewVec_87_T_3[6:0] ? myVec_125 : _GEN_5414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5416 = 7'h7e == _myNewVec_87_T_3[6:0] ? myVec_126 : _GEN_5415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_87 = 7'h7f == _myNewVec_87_T_3[6:0] ? myVec_127 : _GEN_5416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_86_T_3 = _myNewVec_127_T_1 + 16'h29; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_5419 = 7'h1 == _myNewVec_86_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5420 = 7'h2 == _myNewVec_86_T_3[6:0] ? myVec_2 : _GEN_5419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5421 = 7'h3 == _myNewVec_86_T_3[6:0] ? myVec_3 : _GEN_5420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5422 = 7'h4 == _myNewVec_86_T_3[6:0] ? myVec_4 : _GEN_5421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5423 = 7'h5 == _myNewVec_86_T_3[6:0] ? myVec_5 : _GEN_5422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5424 = 7'h6 == _myNewVec_86_T_3[6:0] ? myVec_6 : _GEN_5423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5425 = 7'h7 == _myNewVec_86_T_3[6:0] ? myVec_7 : _GEN_5424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5426 = 7'h8 == _myNewVec_86_T_3[6:0] ? myVec_8 : _GEN_5425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5427 = 7'h9 == _myNewVec_86_T_3[6:0] ? myVec_9 : _GEN_5426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5428 = 7'ha == _myNewVec_86_T_3[6:0] ? myVec_10 : _GEN_5427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5429 = 7'hb == _myNewVec_86_T_3[6:0] ? myVec_11 : _GEN_5428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5430 = 7'hc == _myNewVec_86_T_3[6:0] ? myVec_12 : _GEN_5429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5431 = 7'hd == _myNewVec_86_T_3[6:0] ? myVec_13 : _GEN_5430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5432 = 7'he == _myNewVec_86_T_3[6:0] ? myVec_14 : _GEN_5431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5433 = 7'hf == _myNewVec_86_T_3[6:0] ? myVec_15 : _GEN_5432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5434 = 7'h10 == _myNewVec_86_T_3[6:0] ? myVec_16 : _GEN_5433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5435 = 7'h11 == _myNewVec_86_T_3[6:0] ? myVec_17 : _GEN_5434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5436 = 7'h12 == _myNewVec_86_T_3[6:0] ? myVec_18 : _GEN_5435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5437 = 7'h13 == _myNewVec_86_T_3[6:0] ? myVec_19 : _GEN_5436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5438 = 7'h14 == _myNewVec_86_T_3[6:0] ? myVec_20 : _GEN_5437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5439 = 7'h15 == _myNewVec_86_T_3[6:0] ? myVec_21 : _GEN_5438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5440 = 7'h16 == _myNewVec_86_T_3[6:0] ? myVec_22 : _GEN_5439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5441 = 7'h17 == _myNewVec_86_T_3[6:0] ? myVec_23 : _GEN_5440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5442 = 7'h18 == _myNewVec_86_T_3[6:0] ? myVec_24 : _GEN_5441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5443 = 7'h19 == _myNewVec_86_T_3[6:0] ? myVec_25 : _GEN_5442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5444 = 7'h1a == _myNewVec_86_T_3[6:0] ? myVec_26 : _GEN_5443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5445 = 7'h1b == _myNewVec_86_T_3[6:0] ? myVec_27 : _GEN_5444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5446 = 7'h1c == _myNewVec_86_T_3[6:0] ? myVec_28 : _GEN_5445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5447 = 7'h1d == _myNewVec_86_T_3[6:0] ? myVec_29 : _GEN_5446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5448 = 7'h1e == _myNewVec_86_T_3[6:0] ? myVec_30 : _GEN_5447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5449 = 7'h1f == _myNewVec_86_T_3[6:0] ? myVec_31 : _GEN_5448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5450 = 7'h20 == _myNewVec_86_T_3[6:0] ? myVec_32 : _GEN_5449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5451 = 7'h21 == _myNewVec_86_T_3[6:0] ? myVec_33 : _GEN_5450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5452 = 7'h22 == _myNewVec_86_T_3[6:0] ? myVec_34 : _GEN_5451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5453 = 7'h23 == _myNewVec_86_T_3[6:0] ? myVec_35 : _GEN_5452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5454 = 7'h24 == _myNewVec_86_T_3[6:0] ? myVec_36 : _GEN_5453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5455 = 7'h25 == _myNewVec_86_T_3[6:0] ? myVec_37 : _GEN_5454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5456 = 7'h26 == _myNewVec_86_T_3[6:0] ? myVec_38 : _GEN_5455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5457 = 7'h27 == _myNewVec_86_T_3[6:0] ? myVec_39 : _GEN_5456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5458 = 7'h28 == _myNewVec_86_T_3[6:0] ? myVec_40 : _GEN_5457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5459 = 7'h29 == _myNewVec_86_T_3[6:0] ? myVec_41 : _GEN_5458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5460 = 7'h2a == _myNewVec_86_T_3[6:0] ? myVec_42 : _GEN_5459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5461 = 7'h2b == _myNewVec_86_T_3[6:0] ? myVec_43 : _GEN_5460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5462 = 7'h2c == _myNewVec_86_T_3[6:0] ? myVec_44 : _GEN_5461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5463 = 7'h2d == _myNewVec_86_T_3[6:0] ? myVec_45 : _GEN_5462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5464 = 7'h2e == _myNewVec_86_T_3[6:0] ? myVec_46 : _GEN_5463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5465 = 7'h2f == _myNewVec_86_T_3[6:0] ? myVec_47 : _GEN_5464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5466 = 7'h30 == _myNewVec_86_T_3[6:0] ? myVec_48 : _GEN_5465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5467 = 7'h31 == _myNewVec_86_T_3[6:0] ? myVec_49 : _GEN_5466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5468 = 7'h32 == _myNewVec_86_T_3[6:0] ? myVec_50 : _GEN_5467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5469 = 7'h33 == _myNewVec_86_T_3[6:0] ? myVec_51 : _GEN_5468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5470 = 7'h34 == _myNewVec_86_T_3[6:0] ? myVec_52 : _GEN_5469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5471 = 7'h35 == _myNewVec_86_T_3[6:0] ? myVec_53 : _GEN_5470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5472 = 7'h36 == _myNewVec_86_T_3[6:0] ? myVec_54 : _GEN_5471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5473 = 7'h37 == _myNewVec_86_T_3[6:0] ? myVec_55 : _GEN_5472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5474 = 7'h38 == _myNewVec_86_T_3[6:0] ? myVec_56 : _GEN_5473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5475 = 7'h39 == _myNewVec_86_T_3[6:0] ? myVec_57 : _GEN_5474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5476 = 7'h3a == _myNewVec_86_T_3[6:0] ? myVec_58 : _GEN_5475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5477 = 7'h3b == _myNewVec_86_T_3[6:0] ? myVec_59 : _GEN_5476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5478 = 7'h3c == _myNewVec_86_T_3[6:0] ? myVec_60 : _GEN_5477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5479 = 7'h3d == _myNewVec_86_T_3[6:0] ? myVec_61 : _GEN_5478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5480 = 7'h3e == _myNewVec_86_T_3[6:0] ? myVec_62 : _GEN_5479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5481 = 7'h3f == _myNewVec_86_T_3[6:0] ? myVec_63 : _GEN_5480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5482 = 7'h40 == _myNewVec_86_T_3[6:0] ? myVec_64 : _GEN_5481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5483 = 7'h41 == _myNewVec_86_T_3[6:0] ? myVec_65 : _GEN_5482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5484 = 7'h42 == _myNewVec_86_T_3[6:0] ? myVec_66 : _GEN_5483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5485 = 7'h43 == _myNewVec_86_T_3[6:0] ? myVec_67 : _GEN_5484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5486 = 7'h44 == _myNewVec_86_T_3[6:0] ? myVec_68 : _GEN_5485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5487 = 7'h45 == _myNewVec_86_T_3[6:0] ? myVec_69 : _GEN_5486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5488 = 7'h46 == _myNewVec_86_T_3[6:0] ? myVec_70 : _GEN_5487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5489 = 7'h47 == _myNewVec_86_T_3[6:0] ? myVec_71 : _GEN_5488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5490 = 7'h48 == _myNewVec_86_T_3[6:0] ? myVec_72 : _GEN_5489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5491 = 7'h49 == _myNewVec_86_T_3[6:0] ? myVec_73 : _GEN_5490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5492 = 7'h4a == _myNewVec_86_T_3[6:0] ? myVec_74 : _GEN_5491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5493 = 7'h4b == _myNewVec_86_T_3[6:0] ? myVec_75 : _GEN_5492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5494 = 7'h4c == _myNewVec_86_T_3[6:0] ? myVec_76 : _GEN_5493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5495 = 7'h4d == _myNewVec_86_T_3[6:0] ? myVec_77 : _GEN_5494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5496 = 7'h4e == _myNewVec_86_T_3[6:0] ? myVec_78 : _GEN_5495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5497 = 7'h4f == _myNewVec_86_T_3[6:0] ? myVec_79 : _GEN_5496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5498 = 7'h50 == _myNewVec_86_T_3[6:0] ? myVec_80 : _GEN_5497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5499 = 7'h51 == _myNewVec_86_T_3[6:0] ? myVec_81 : _GEN_5498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5500 = 7'h52 == _myNewVec_86_T_3[6:0] ? myVec_82 : _GEN_5499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5501 = 7'h53 == _myNewVec_86_T_3[6:0] ? myVec_83 : _GEN_5500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5502 = 7'h54 == _myNewVec_86_T_3[6:0] ? myVec_84 : _GEN_5501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5503 = 7'h55 == _myNewVec_86_T_3[6:0] ? myVec_85 : _GEN_5502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5504 = 7'h56 == _myNewVec_86_T_3[6:0] ? myVec_86 : _GEN_5503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5505 = 7'h57 == _myNewVec_86_T_3[6:0] ? myVec_87 : _GEN_5504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5506 = 7'h58 == _myNewVec_86_T_3[6:0] ? myVec_88 : _GEN_5505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5507 = 7'h59 == _myNewVec_86_T_3[6:0] ? myVec_89 : _GEN_5506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5508 = 7'h5a == _myNewVec_86_T_3[6:0] ? myVec_90 : _GEN_5507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5509 = 7'h5b == _myNewVec_86_T_3[6:0] ? myVec_91 : _GEN_5508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5510 = 7'h5c == _myNewVec_86_T_3[6:0] ? myVec_92 : _GEN_5509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5511 = 7'h5d == _myNewVec_86_T_3[6:0] ? myVec_93 : _GEN_5510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5512 = 7'h5e == _myNewVec_86_T_3[6:0] ? myVec_94 : _GEN_5511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5513 = 7'h5f == _myNewVec_86_T_3[6:0] ? myVec_95 : _GEN_5512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5514 = 7'h60 == _myNewVec_86_T_3[6:0] ? myVec_96 : _GEN_5513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5515 = 7'h61 == _myNewVec_86_T_3[6:0] ? myVec_97 : _GEN_5514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5516 = 7'h62 == _myNewVec_86_T_3[6:0] ? myVec_98 : _GEN_5515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5517 = 7'h63 == _myNewVec_86_T_3[6:0] ? myVec_99 : _GEN_5516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5518 = 7'h64 == _myNewVec_86_T_3[6:0] ? myVec_100 : _GEN_5517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5519 = 7'h65 == _myNewVec_86_T_3[6:0] ? myVec_101 : _GEN_5518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5520 = 7'h66 == _myNewVec_86_T_3[6:0] ? myVec_102 : _GEN_5519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5521 = 7'h67 == _myNewVec_86_T_3[6:0] ? myVec_103 : _GEN_5520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5522 = 7'h68 == _myNewVec_86_T_3[6:0] ? myVec_104 : _GEN_5521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5523 = 7'h69 == _myNewVec_86_T_3[6:0] ? myVec_105 : _GEN_5522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5524 = 7'h6a == _myNewVec_86_T_3[6:0] ? myVec_106 : _GEN_5523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5525 = 7'h6b == _myNewVec_86_T_3[6:0] ? myVec_107 : _GEN_5524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5526 = 7'h6c == _myNewVec_86_T_3[6:0] ? myVec_108 : _GEN_5525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5527 = 7'h6d == _myNewVec_86_T_3[6:0] ? myVec_109 : _GEN_5526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5528 = 7'h6e == _myNewVec_86_T_3[6:0] ? myVec_110 : _GEN_5527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5529 = 7'h6f == _myNewVec_86_T_3[6:0] ? myVec_111 : _GEN_5528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5530 = 7'h70 == _myNewVec_86_T_3[6:0] ? myVec_112 : _GEN_5529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5531 = 7'h71 == _myNewVec_86_T_3[6:0] ? myVec_113 : _GEN_5530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5532 = 7'h72 == _myNewVec_86_T_3[6:0] ? myVec_114 : _GEN_5531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5533 = 7'h73 == _myNewVec_86_T_3[6:0] ? myVec_115 : _GEN_5532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5534 = 7'h74 == _myNewVec_86_T_3[6:0] ? myVec_116 : _GEN_5533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5535 = 7'h75 == _myNewVec_86_T_3[6:0] ? myVec_117 : _GEN_5534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5536 = 7'h76 == _myNewVec_86_T_3[6:0] ? myVec_118 : _GEN_5535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5537 = 7'h77 == _myNewVec_86_T_3[6:0] ? myVec_119 : _GEN_5536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5538 = 7'h78 == _myNewVec_86_T_3[6:0] ? myVec_120 : _GEN_5537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5539 = 7'h79 == _myNewVec_86_T_3[6:0] ? myVec_121 : _GEN_5538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5540 = 7'h7a == _myNewVec_86_T_3[6:0] ? myVec_122 : _GEN_5539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5541 = 7'h7b == _myNewVec_86_T_3[6:0] ? myVec_123 : _GEN_5540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5542 = 7'h7c == _myNewVec_86_T_3[6:0] ? myVec_124 : _GEN_5541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5543 = 7'h7d == _myNewVec_86_T_3[6:0] ? myVec_125 : _GEN_5542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5544 = 7'h7e == _myNewVec_86_T_3[6:0] ? myVec_126 : _GEN_5543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_86 = 7'h7f == _myNewVec_86_T_3[6:0] ? myVec_127 : _GEN_5544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_85_T_3 = _myNewVec_127_T_1 + 16'h2a; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_5547 = 7'h1 == _myNewVec_85_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5548 = 7'h2 == _myNewVec_85_T_3[6:0] ? myVec_2 : _GEN_5547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5549 = 7'h3 == _myNewVec_85_T_3[6:0] ? myVec_3 : _GEN_5548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5550 = 7'h4 == _myNewVec_85_T_3[6:0] ? myVec_4 : _GEN_5549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5551 = 7'h5 == _myNewVec_85_T_3[6:0] ? myVec_5 : _GEN_5550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5552 = 7'h6 == _myNewVec_85_T_3[6:0] ? myVec_6 : _GEN_5551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5553 = 7'h7 == _myNewVec_85_T_3[6:0] ? myVec_7 : _GEN_5552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5554 = 7'h8 == _myNewVec_85_T_3[6:0] ? myVec_8 : _GEN_5553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5555 = 7'h9 == _myNewVec_85_T_3[6:0] ? myVec_9 : _GEN_5554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5556 = 7'ha == _myNewVec_85_T_3[6:0] ? myVec_10 : _GEN_5555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5557 = 7'hb == _myNewVec_85_T_3[6:0] ? myVec_11 : _GEN_5556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5558 = 7'hc == _myNewVec_85_T_3[6:0] ? myVec_12 : _GEN_5557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5559 = 7'hd == _myNewVec_85_T_3[6:0] ? myVec_13 : _GEN_5558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5560 = 7'he == _myNewVec_85_T_3[6:0] ? myVec_14 : _GEN_5559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5561 = 7'hf == _myNewVec_85_T_3[6:0] ? myVec_15 : _GEN_5560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5562 = 7'h10 == _myNewVec_85_T_3[6:0] ? myVec_16 : _GEN_5561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5563 = 7'h11 == _myNewVec_85_T_3[6:0] ? myVec_17 : _GEN_5562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5564 = 7'h12 == _myNewVec_85_T_3[6:0] ? myVec_18 : _GEN_5563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5565 = 7'h13 == _myNewVec_85_T_3[6:0] ? myVec_19 : _GEN_5564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5566 = 7'h14 == _myNewVec_85_T_3[6:0] ? myVec_20 : _GEN_5565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5567 = 7'h15 == _myNewVec_85_T_3[6:0] ? myVec_21 : _GEN_5566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5568 = 7'h16 == _myNewVec_85_T_3[6:0] ? myVec_22 : _GEN_5567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5569 = 7'h17 == _myNewVec_85_T_3[6:0] ? myVec_23 : _GEN_5568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5570 = 7'h18 == _myNewVec_85_T_3[6:0] ? myVec_24 : _GEN_5569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5571 = 7'h19 == _myNewVec_85_T_3[6:0] ? myVec_25 : _GEN_5570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5572 = 7'h1a == _myNewVec_85_T_3[6:0] ? myVec_26 : _GEN_5571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5573 = 7'h1b == _myNewVec_85_T_3[6:0] ? myVec_27 : _GEN_5572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5574 = 7'h1c == _myNewVec_85_T_3[6:0] ? myVec_28 : _GEN_5573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5575 = 7'h1d == _myNewVec_85_T_3[6:0] ? myVec_29 : _GEN_5574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5576 = 7'h1e == _myNewVec_85_T_3[6:0] ? myVec_30 : _GEN_5575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5577 = 7'h1f == _myNewVec_85_T_3[6:0] ? myVec_31 : _GEN_5576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5578 = 7'h20 == _myNewVec_85_T_3[6:0] ? myVec_32 : _GEN_5577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5579 = 7'h21 == _myNewVec_85_T_3[6:0] ? myVec_33 : _GEN_5578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5580 = 7'h22 == _myNewVec_85_T_3[6:0] ? myVec_34 : _GEN_5579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5581 = 7'h23 == _myNewVec_85_T_3[6:0] ? myVec_35 : _GEN_5580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5582 = 7'h24 == _myNewVec_85_T_3[6:0] ? myVec_36 : _GEN_5581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5583 = 7'h25 == _myNewVec_85_T_3[6:0] ? myVec_37 : _GEN_5582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5584 = 7'h26 == _myNewVec_85_T_3[6:0] ? myVec_38 : _GEN_5583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5585 = 7'h27 == _myNewVec_85_T_3[6:0] ? myVec_39 : _GEN_5584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5586 = 7'h28 == _myNewVec_85_T_3[6:0] ? myVec_40 : _GEN_5585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5587 = 7'h29 == _myNewVec_85_T_3[6:0] ? myVec_41 : _GEN_5586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5588 = 7'h2a == _myNewVec_85_T_3[6:0] ? myVec_42 : _GEN_5587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5589 = 7'h2b == _myNewVec_85_T_3[6:0] ? myVec_43 : _GEN_5588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5590 = 7'h2c == _myNewVec_85_T_3[6:0] ? myVec_44 : _GEN_5589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5591 = 7'h2d == _myNewVec_85_T_3[6:0] ? myVec_45 : _GEN_5590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5592 = 7'h2e == _myNewVec_85_T_3[6:0] ? myVec_46 : _GEN_5591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5593 = 7'h2f == _myNewVec_85_T_3[6:0] ? myVec_47 : _GEN_5592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5594 = 7'h30 == _myNewVec_85_T_3[6:0] ? myVec_48 : _GEN_5593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5595 = 7'h31 == _myNewVec_85_T_3[6:0] ? myVec_49 : _GEN_5594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5596 = 7'h32 == _myNewVec_85_T_3[6:0] ? myVec_50 : _GEN_5595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5597 = 7'h33 == _myNewVec_85_T_3[6:0] ? myVec_51 : _GEN_5596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5598 = 7'h34 == _myNewVec_85_T_3[6:0] ? myVec_52 : _GEN_5597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5599 = 7'h35 == _myNewVec_85_T_3[6:0] ? myVec_53 : _GEN_5598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5600 = 7'h36 == _myNewVec_85_T_3[6:0] ? myVec_54 : _GEN_5599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5601 = 7'h37 == _myNewVec_85_T_3[6:0] ? myVec_55 : _GEN_5600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5602 = 7'h38 == _myNewVec_85_T_3[6:0] ? myVec_56 : _GEN_5601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5603 = 7'h39 == _myNewVec_85_T_3[6:0] ? myVec_57 : _GEN_5602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5604 = 7'h3a == _myNewVec_85_T_3[6:0] ? myVec_58 : _GEN_5603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5605 = 7'h3b == _myNewVec_85_T_3[6:0] ? myVec_59 : _GEN_5604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5606 = 7'h3c == _myNewVec_85_T_3[6:0] ? myVec_60 : _GEN_5605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5607 = 7'h3d == _myNewVec_85_T_3[6:0] ? myVec_61 : _GEN_5606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5608 = 7'h3e == _myNewVec_85_T_3[6:0] ? myVec_62 : _GEN_5607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5609 = 7'h3f == _myNewVec_85_T_3[6:0] ? myVec_63 : _GEN_5608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5610 = 7'h40 == _myNewVec_85_T_3[6:0] ? myVec_64 : _GEN_5609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5611 = 7'h41 == _myNewVec_85_T_3[6:0] ? myVec_65 : _GEN_5610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5612 = 7'h42 == _myNewVec_85_T_3[6:0] ? myVec_66 : _GEN_5611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5613 = 7'h43 == _myNewVec_85_T_3[6:0] ? myVec_67 : _GEN_5612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5614 = 7'h44 == _myNewVec_85_T_3[6:0] ? myVec_68 : _GEN_5613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5615 = 7'h45 == _myNewVec_85_T_3[6:0] ? myVec_69 : _GEN_5614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5616 = 7'h46 == _myNewVec_85_T_3[6:0] ? myVec_70 : _GEN_5615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5617 = 7'h47 == _myNewVec_85_T_3[6:0] ? myVec_71 : _GEN_5616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5618 = 7'h48 == _myNewVec_85_T_3[6:0] ? myVec_72 : _GEN_5617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5619 = 7'h49 == _myNewVec_85_T_3[6:0] ? myVec_73 : _GEN_5618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5620 = 7'h4a == _myNewVec_85_T_3[6:0] ? myVec_74 : _GEN_5619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5621 = 7'h4b == _myNewVec_85_T_3[6:0] ? myVec_75 : _GEN_5620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5622 = 7'h4c == _myNewVec_85_T_3[6:0] ? myVec_76 : _GEN_5621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5623 = 7'h4d == _myNewVec_85_T_3[6:0] ? myVec_77 : _GEN_5622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5624 = 7'h4e == _myNewVec_85_T_3[6:0] ? myVec_78 : _GEN_5623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5625 = 7'h4f == _myNewVec_85_T_3[6:0] ? myVec_79 : _GEN_5624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5626 = 7'h50 == _myNewVec_85_T_3[6:0] ? myVec_80 : _GEN_5625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5627 = 7'h51 == _myNewVec_85_T_3[6:0] ? myVec_81 : _GEN_5626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5628 = 7'h52 == _myNewVec_85_T_3[6:0] ? myVec_82 : _GEN_5627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5629 = 7'h53 == _myNewVec_85_T_3[6:0] ? myVec_83 : _GEN_5628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5630 = 7'h54 == _myNewVec_85_T_3[6:0] ? myVec_84 : _GEN_5629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5631 = 7'h55 == _myNewVec_85_T_3[6:0] ? myVec_85 : _GEN_5630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5632 = 7'h56 == _myNewVec_85_T_3[6:0] ? myVec_86 : _GEN_5631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5633 = 7'h57 == _myNewVec_85_T_3[6:0] ? myVec_87 : _GEN_5632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5634 = 7'h58 == _myNewVec_85_T_3[6:0] ? myVec_88 : _GEN_5633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5635 = 7'h59 == _myNewVec_85_T_3[6:0] ? myVec_89 : _GEN_5634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5636 = 7'h5a == _myNewVec_85_T_3[6:0] ? myVec_90 : _GEN_5635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5637 = 7'h5b == _myNewVec_85_T_3[6:0] ? myVec_91 : _GEN_5636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5638 = 7'h5c == _myNewVec_85_T_3[6:0] ? myVec_92 : _GEN_5637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5639 = 7'h5d == _myNewVec_85_T_3[6:0] ? myVec_93 : _GEN_5638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5640 = 7'h5e == _myNewVec_85_T_3[6:0] ? myVec_94 : _GEN_5639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5641 = 7'h5f == _myNewVec_85_T_3[6:0] ? myVec_95 : _GEN_5640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5642 = 7'h60 == _myNewVec_85_T_3[6:0] ? myVec_96 : _GEN_5641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5643 = 7'h61 == _myNewVec_85_T_3[6:0] ? myVec_97 : _GEN_5642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5644 = 7'h62 == _myNewVec_85_T_3[6:0] ? myVec_98 : _GEN_5643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5645 = 7'h63 == _myNewVec_85_T_3[6:0] ? myVec_99 : _GEN_5644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5646 = 7'h64 == _myNewVec_85_T_3[6:0] ? myVec_100 : _GEN_5645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5647 = 7'h65 == _myNewVec_85_T_3[6:0] ? myVec_101 : _GEN_5646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5648 = 7'h66 == _myNewVec_85_T_3[6:0] ? myVec_102 : _GEN_5647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5649 = 7'h67 == _myNewVec_85_T_3[6:0] ? myVec_103 : _GEN_5648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5650 = 7'h68 == _myNewVec_85_T_3[6:0] ? myVec_104 : _GEN_5649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5651 = 7'h69 == _myNewVec_85_T_3[6:0] ? myVec_105 : _GEN_5650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5652 = 7'h6a == _myNewVec_85_T_3[6:0] ? myVec_106 : _GEN_5651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5653 = 7'h6b == _myNewVec_85_T_3[6:0] ? myVec_107 : _GEN_5652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5654 = 7'h6c == _myNewVec_85_T_3[6:0] ? myVec_108 : _GEN_5653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5655 = 7'h6d == _myNewVec_85_T_3[6:0] ? myVec_109 : _GEN_5654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5656 = 7'h6e == _myNewVec_85_T_3[6:0] ? myVec_110 : _GEN_5655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5657 = 7'h6f == _myNewVec_85_T_3[6:0] ? myVec_111 : _GEN_5656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5658 = 7'h70 == _myNewVec_85_T_3[6:0] ? myVec_112 : _GEN_5657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5659 = 7'h71 == _myNewVec_85_T_3[6:0] ? myVec_113 : _GEN_5658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5660 = 7'h72 == _myNewVec_85_T_3[6:0] ? myVec_114 : _GEN_5659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5661 = 7'h73 == _myNewVec_85_T_3[6:0] ? myVec_115 : _GEN_5660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5662 = 7'h74 == _myNewVec_85_T_3[6:0] ? myVec_116 : _GEN_5661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5663 = 7'h75 == _myNewVec_85_T_3[6:0] ? myVec_117 : _GEN_5662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5664 = 7'h76 == _myNewVec_85_T_3[6:0] ? myVec_118 : _GEN_5663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5665 = 7'h77 == _myNewVec_85_T_3[6:0] ? myVec_119 : _GEN_5664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5666 = 7'h78 == _myNewVec_85_T_3[6:0] ? myVec_120 : _GEN_5665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5667 = 7'h79 == _myNewVec_85_T_3[6:0] ? myVec_121 : _GEN_5666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5668 = 7'h7a == _myNewVec_85_T_3[6:0] ? myVec_122 : _GEN_5667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5669 = 7'h7b == _myNewVec_85_T_3[6:0] ? myVec_123 : _GEN_5668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5670 = 7'h7c == _myNewVec_85_T_3[6:0] ? myVec_124 : _GEN_5669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5671 = 7'h7d == _myNewVec_85_T_3[6:0] ? myVec_125 : _GEN_5670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5672 = 7'h7e == _myNewVec_85_T_3[6:0] ? myVec_126 : _GEN_5671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_85 = 7'h7f == _myNewVec_85_T_3[6:0] ? myVec_127 : _GEN_5672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_84_T_3 = _myNewVec_127_T_1 + 16'h2b; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_5675 = 7'h1 == _myNewVec_84_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5676 = 7'h2 == _myNewVec_84_T_3[6:0] ? myVec_2 : _GEN_5675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5677 = 7'h3 == _myNewVec_84_T_3[6:0] ? myVec_3 : _GEN_5676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5678 = 7'h4 == _myNewVec_84_T_3[6:0] ? myVec_4 : _GEN_5677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5679 = 7'h5 == _myNewVec_84_T_3[6:0] ? myVec_5 : _GEN_5678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5680 = 7'h6 == _myNewVec_84_T_3[6:0] ? myVec_6 : _GEN_5679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5681 = 7'h7 == _myNewVec_84_T_3[6:0] ? myVec_7 : _GEN_5680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5682 = 7'h8 == _myNewVec_84_T_3[6:0] ? myVec_8 : _GEN_5681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5683 = 7'h9 == _myNewVec_84_T_3[6:0] ? myVec_9 : _GEN_5682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5684 = 7'ha == _myNewVec_84_T_3[6:0] ? myVec_10 : _GEN_5683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5685 = 7'hb == _myNewVec_84_T_3[6:0] ? myVec_11 : _GEN_5684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5686 = 7'hc == _myNewVec_84_T_3[6:0] ? myVec_12 : _GEN_5685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5687 = 7'hd == _myNewVec_84_T_3[6:0] ? myVec_13 : _GEN_5686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5688 = 7'he == _myNewVec_84_T_3[6:0] ? myVec_14 : _GEN_5687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5689 = 7'hf == _myNewVec_84_T_3[6:0] ? myVec_15 : _GEN_5688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5690 = 7'h10 == _myNewVec_84_T_3[6:0] ? myVec_16 : _GEN_5689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5691 = 7'h11 == _myNewVec_84_T_3[6:0] ? myVec_17 : _GEN_5690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5692 = 7'h12 == _myNewVec_84_T_3[6:0] ? myVec_18 : _GEN_5691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5693 = 7'h13 == _myNewVec_84_T_3[6:0] ? myVec_19 : _GEN_5692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5694 = 7'h14 == _myNewVec_84_T_3[6:0] ? myVec_20 : _GEN_5693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5695 = 7'h15 == _myNewVec_84_T_3[6:0] ? myVec_21 : _GEN_5694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5696 = 7'h16 == _myNewVec_84_T_3[6:0] ? myVec_22 : _GEN_5695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5697 = 7'h17 == _myNewVec_84_T_3[6:0] ? myVec_23 : _GEN_5696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5698 = 7'h18 == _myNewVec_84_T_3[6:0] ? myVec_24 : _GEN_5697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5699 = 7'h19 == _myNewVec_84_T_3[6:0] ? myVec_25 : _GEN_5698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5700 = 7'h1a == _myNewVec_84_T_3[6:0] ? myVec_26 : _GEN_5699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5701 = 7'h1b == _myNewVec_84_T_3[6:0] ? myVec_27 : _GEN_5700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5702 = 7'h1c == _myNewVec_84_T_3[6:0] ? myVec_28 : _GEN_5701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5703 = 7'h1d == _myNewVec_84_T_3[6:0] ? myVec_29 : _GEN_5702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5704 = 7'h1e == _myNewVec_84_T_3[6:0] ? myVec_30 : _GEN_5703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5705 = 7'h1f == _myNewVec_84_T_3[6:0] ? myVec_31 : _GEN_5704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5706 = 7'h20 == _myNewVec_84_T_3[6:0] ? myVec_32 : _GEN_5705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5707 = 7'h21 == _myNewVec_84_T_3[6:0] ? myVec_33 : _GEN_5706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5708 = 7'h22 == _myNewVec_84_T_3[6:0] ? myVec_34 : _GEN_5707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5709 = 7'h23 == _myNewVec_84_T_3[6:0] ? myVec_35 : _GEN_5708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5710 = 7'h24 == _myNewVec_84_T_3[6:0] ? myVec_36 : _GEN_5709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5711 = 7'h25 == _myNewVec_84_T_3[6:0] ? myVec_37 : _GEN_5710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5712 = 7'h26 == _myNewVec_84_T_3[6:0] ? myVec_38 : _GEN_5711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5713 = 7'h27 == _myNewVec_84_T_3[6:0] ? myVec_39 : _GEN_5712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5714 = 7'h28 == _myNewVec_84_T_3[6:0] ? myVec_40 : _GEN_5713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5715 = 7'h29 == _myNewVec_84_T_3[6:0] ? myVec_41 : _GEN_5714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5716 = 7'h2a == _myNewVec_84_T_3[6:0] ? myVec_42 : _GEN_5715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5717 = 7'h2b == _myNewVec_84_T_3[6:0] ? myVec_43 : _GEN_5716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5718 = 7'h2c == _myNewVec_84_T_3[6:0] ? myVec_44 : _GEN_5717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5719 = 7'h2d == _myNewVec_84_T_3[6:0] ? myVec_45 : _GEN_5718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5720 = 7'h2e == _myNewVec_84_T_3[6:0] ? myVec_46 : _GEN_5719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5721 = 7'h2f == _myNewVec_84_T_3[6:0] ? myVec_47 : _GEN_5720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5722 = 7'h30 == _myNewVec_84_T_3[6:0] ? myVec_48 : _GEN_5721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5723 = 7'h31 == _myNewVec_84_T_3[6:0] ? myVec_49 : _GEN_5722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5724 = 7'h32 == _myNewVec_84_T_3[6:0] ? myVec_50 : _GEN_5723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5725 = 7'h33 == _myNewVec_84_T_3[6:0] ? myVec_51 : _GEN_5724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5726 = 7'h34 == _myNewVec_84_T_3[6:0] ? myVec_52 : _GEN_5725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5727 = 7'h35 == _myNewVec_84_T_3[6:0] ? myVec_53 : _GEN_5726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5728 = 7'h36 == _myNewVec_84_T_3[6:0] ? myVec_54 : _GEN_5727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5729 = 7'h37 == _myNewVec_84_T_3[6:0] ? myVec_55 : _GEN_5728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5730 = 7'h38 == _myNewVec_84_T_3[6:0] ? myVec_56 : _GEN_5729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5731 = 7'h39 == _myNewVec_84_T_3[6:0] ? myVec_57 : _GEN_5730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5732 = 7'h3a == _myNewVec_84_T_3[6:0] ? myVec_58 : _GEN_5731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5733 = 7'h3b == _myNewVec_84_T_3[6:0] ? myVec_59 : _GEN_5732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5734 = 7'h3c == _myNewVec_84_T_3[6:0] ? myVec_60 : _GEN_5733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5735 = 7'h3d == _myNewVec_84_T_3[6:0] ? myVec_61 : _GEN_5734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5736 = 7'h3e == _myNewVec_84_T_3[6:0] ? myVec_62 : _GEN_5735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5737 = 7'h3f == _myNewVec_84_T_3[6:0] ? myVec_63 : _GEN_5736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5738 = 7'h40 == _myNewVec_84_T_3[6:0] ? myVec_64 : _GEN_5737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5739 = 7'h41 == _myNewVec_84_T_3[6:0] ? myVec_65 : _GEN_5738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5740 = 7'h42 == _myNewVec_84_T_3[6:0] ? myVec_66 : _GEN_5739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5741 = 7'h43 == _myNewVec_84_T_3[6:0] ? myVec_67 : _GEN_5740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5742 = 7'h44 == _myNewVec_84_T_3[6:0] ? myVec_68 : _GEN_5741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5743 = 7'h45 == _myNewVec_84_T_3[6:0] ? myVec_69 : _GEN_5742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5744 = 7'h46 == _myNewVec_84_T_3[6:0] ? myVec_70 : _GEN_5743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5745 = 7'h47 == _myNewVec_84_T_3[6:0] ? myVec_71 : _GEN_5744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5746 = 7'h48 == _myNewVec_84_T_3[6:0] ? myVec_72 : _GEN_5745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5747 = 7'h49 == _myNewVec_84_T_3[6:0] ? myVec_73 : _GEN_5746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5748 = 7'h4a == _myNewVec_84_T_3[6:0] ? myVec_74 : _GEN_5747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5749 = 7'h4b == _myNewVec_84_T_3[6:0] ? myVec_75 : _GEN_5748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5750 = 7'h4c == _myNewVec_84_T_3[6:0] ? myVec_76 : _GEN_5749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5751 = 7'h4d == _myNewVec_84_T_3[6:0] ? myVec_77 : _GEN_5750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5752 = 7'h4e == _myNewVec_84_T_3[6:0] ? myVec_78 : _GEN_5751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5753 = 7'h4f == _myNewVec_84_T_3[6:0] ? myVec_79 : _GEN_5752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5754 = 7'h50 == _myNewVec_84_T_3[6:0] ? myVec_80 : _GEN_5753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5755 = 7'h51 == _myNewVec_84_T_3[6:0] ? myVec_81 : _GEN_5754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5756 = 7'h52 == _myNewVec_84_T_3[6:0] ? myVec_82 : _GEN_5755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5757 = 7'h53 == _myNewVec_84_T_3[6:0] ? myVec_83 : _GEN_5756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5758 = 7'h54 == _myNewVec_84_T_3[6:0] ? myVec_84 : _GEN_5757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5759 = 7'h55 == _myNewVec_84_T_3[6:0] ? myVec_85 : _GEN_5758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5760 = 7'h56 == _myNewVec_84_T_3[6:0] ? myVec_86 : _GEN_5759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5761 = 7'h57 == _myNewVec_84_T_3[6:0] ? myVec_87 : _GEN_5760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5762 = 7'h58 == _myNewVec_84_T_3[6:0] ? myVec_88 : _GEN_5761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5763 = 7'h59 == _myNewVec_84_T_3[6:0] ? myVec_89 : _GEN_5762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5764 = 7'h5a == _myNewVec_84_T_3[6:0] ? myVec_90 : _GEN_5763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5765 = 7'h5b == _myNewVec_84_T_3[6:0] ? myVec_91 : _GEN_5764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5766 = 7'h5c == _myNewVec_84_T_3[6:0] ? myVec_92 : _GEN_5765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5767 = 7'h5d == _myNewVec_84_T_3[6:0] ? myVec_93 : _GEN_5766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5768 = 7'h5e == _myNewVec_84_T_3[6:0] ? myVec_94 : _GEN_5767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5769 = 7'h5f == _myNewVec_84_T_3[6:0] ? myVec_95 : _GEN_5768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5770 = 7'h60 == _myNewVec_84_T_3[6:0] ? myVec_96 : _GEN_5769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5771 = 7'h61 == _myNewVec_84_T_3[6:0] ? myVec_97 : _GEN_5770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5772 = 7'h62 == _myNewVec_84_T_3[6:0] ? myVec_98 : _GEN_5771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5773 = 7'h63 == _myNewVec_84_T_3[6:0] ? myVec_99 : _GEN_5772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5774 = 7'h64 == _myNewVec_84_T_3[6:0] ? myVec_100 : _GEN_5773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5775 = 7'h65 == _myNewVec_84_T_3[6:0] ? myVec_101 : _GEN_5774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5776 = 7'h66 == _myNewVec_84_T_3[6:0] ? myVec_102 : _GEN_5775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5777 = 7'h67 == _myNewVec_84_T_3[6:0] ? myVec_103 : _GEN_5776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5778 = 7'h68 == _myNewVec_84_T_3[6:0] ? myVec_104 : _GEN_5777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5779 = 7'h69 == _myNewVec_84_T_3[6:0] ? myVec_105 : _GEN_5778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5780 = 7'h6a == _myNewVec_84_T_3[6:0] ? myVec_106 : _GEN_5779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5781 = 7'h6b == _myNewVec_84_T_3[6:0] ? myVec_107 : _GEN_5780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5782 = 7'h6c == _myNewVec_84_T_3[6:0] ? myVec_108 : _GEN_5781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5783 = 7'h6d == _myNewVec_84_T_3[6:0] ? myVec_109 : _GEN_5782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5784 = 7'h6e == _myNewVec_84_T_3[6:0] ? myVec_110 : _GEN_5783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5785 = 7'h6f == _myNewVec_84_T_3[6:0] ? myVec_111 : _GEN_5784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5786 = 7'h70 == _myNewVec_84_T_3[6:0] ? myVec_112 : _GEN_5785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5787 = 7'h71 == _myNewVec_84_T_3[6:0] ? myVec_113 : _GEN_5786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5788 = 7'h72 == _myNewVec_84_T_3[6:0] ? myVec_114 : _GEN_5787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5789 = 7'h73 == _myNewVec_84_T_3[6:0] ? myVec_115 : _GEN_5788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5790 = 7'h74 == _myNewVec_84_T_3[6:0] ? myVec_116 : _GEN_5789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5791 = 7'h75 == _myNewVec_84_T_3[6:0] ? myVec_117 : _GEN_5790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5792 = 7'h76 == _myNewVec_84_T_3[6:0] ? myVec_118 : _GEN_5791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5793 = 7'h77 == _myNewVec_84_T_3[6:0] ? myVec_119 : _GEN_5792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5794 = 7'h78 == _myNewVec_84_T_3[6:0] ? myVec_120 : _GEN_5793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5795 = 7'h79 == _myNewVec_84_T_3[6:0] ? myVec_121 : _GEN_5794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5796 = 7'h7a == _myNewVec_84_T_3[6:0] ? myVec_122 : _GEN_5795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5797 = 7'h7b == _myNewVec_84_T_3[6:0] ? myVec_123 : _GEN_5796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5798 = 7'h7c == _myNewVec_84_T_3[6:0] ? myVec_124 : _GEN_5797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5799 = 7'h7d == _myNewVec_84_T_3[6:0] ? myVec_125 : _GEN_5798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5800 = 7'h7e == _myNewVec_84_T_3[6:0] ? myVec_126 : _GEN_5799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_84 = 7'h7f == _myNewVec_84_T_3[6:0] ? myVec_127 : _GEN_5800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_83_T_3 = _myNewVec_127_T_1 + 16'h2c; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_5803 = 7'h1 == _myNewVec_83_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5804 = 7'h2 == _myNewVec_83_T_3[6:0] ? myVec_2 : _GEN_5803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5805 = 7'h3 == _myNewVec_83_T_3[6:0] ? myVec_3 : _GEN_5804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5806 = 7'h4 == _myNewVec_83_T_3[6:0] ? myVec_4 : _GEN_5805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5807 = 7'h5 == _myNewVec_83_T_3[6:0] ? myVec_5 : _GEN_5806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5808 = 7'h6 == _myNewVec_83_T_3[6:0] ? myVec_6 : _GEN_5807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5809 = 7'h7 == _myNewVec_83_T_3[6:0] ? myVec_7 : _GEN_5808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5810 = 7'h8 == _myNewVec_83_T_3[6:0] ? myVec_8 : _GEN_5809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5811 = 7'h9 == _myNewVec_83_T_3[6:0] ? myVec_9 : _GEN_5810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5812 = 7'ha == _myNewVec_83_T_3[6:0] ? myVec_10 : _GEN_5811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5813 = 7'hb == _myNewVec_83_T_3[6:0] ? myVec_11 : _GEN_5812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5814 = 7'hc == _myNewVec_83_T_3[6:0] ? myVec_12 : _GEN_5813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5815 = 7'hd == _myNewVec_83_T_3[6:0] ? myVec_13 : _GEN_5814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5816 = 7'he == _myNewVec_83_T_3[6:0] ? myVec_14 : _GEN_5815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5817 = 7'hf == _myNewVec_83_T_3[6:0] ? myVec_15 : _GEN_5816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5818 = 7'h10 == _myNewVec_83_T_3[6:0] ? myVec_16 : _GEN_5817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5819 = 7'h11 == _myNewVec_83_T_3[6:0] ? myVec_17 : _GEN_5818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5820 = 7'h12 == _myNewVec_83_T_3[6:0] ? myVec_18 : _GEN_5819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5821 = 7'h13 == _myNewVec_83_T_3[6:0] ? myVec_19 : _GEN_5820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5822 = 7'h14 == _myNewVec_83_T_3[6:0] ? myVec_20 : _GEN_5821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5823 = 7'h15 == _myNewVec_83_T_3[6:0] ? myVec_21 : _GEN_5822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5824 = 7'h16 == _myNewVec_83_T_3[6:0] ? myVec_22 : _GEN_5823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5825 = 7'h17 == _myNewVec_83_T_3[6:0] ? myVec_23 : _GEN_5824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5826 = 7'h18 == _myNewVec_83_T_3[6:0] ? myVec_24 : _GEN_5825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5827 = 7'h19 == _myNewVec_83_T_3[6:0] ? myVec_25 : _GEN_5826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5828 = 7'h1a == _myNewVec_83_T_3[6:0] ? myVec_26 : _GEN_5827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5829 = 7'h1b == _myNewVec_83_T_3[6:0] ? myVec_27 : _GEN_5828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5830 = 7'h1c == _myNewVec_83_T_3[6:0] ? myVec_28 : _GEN_5829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5831 = 7'h1d == _myNewVec_83_T_3[6:0] ? myVec_29 : _GEN_5830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5832 = 7'h1e == _myNewVec_83_T_3[6:0] ? myVec_30 : _GEN_5831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5833 = 7'h1f == _myNewVec_83_T_3[6:0] ? myVec_31 : _GEN_5832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5834 = 7'h20 == _myNewVec_83_T_3[6:0] ? myVec_32 : _GEN_5833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5835 = 7'h21 == _myNewVec_83_T_3[6:0] ? myVec_33 : _GEN_5834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5836 = 7'h22 == _myNewVec_83_T_3[6:0] ? myVec_34 : _GEN_5835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5837 = 7'h23 == _myNewVec_83_T_3[6:0] ? myVec_35 : _GEN_5836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5838 = 7'h24 == _myNewVec_83_T_3[6:0] ? myVec_36 : _GEN_5837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5839 = 7'h25 == _myNewVec_83_T_3[6:0] ? myVec_37 : _GEN_5838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5840 = 7'h26 == _myNewVec_83_T_3[6:0] ? myVec_38 : _GEN_5839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5841 = 7'h27 == _myNewVec_83_T_3[6:0] ? myVec_39 : _GEN_5840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5842 = 7'h28 == _myNewVec_83_T_3[6:0] ? myVec_40 : _GEN_5841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5843 = 7'h29 == _myNewVec_83_T_3[6:0] ? myVec_41 : _GEN_5842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5844 = 7'h2a == _myNewVec_83_T_3[6:0] ? myVec_42 : _GEN_5843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5845 = 7'h2b == _myNewVec_83_T_3[6:0] ? myVec_43 : _GEN_5844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5846 = 7'h2c == _myNewVec_83_T_3[6:0] ? myVec_44 : _GEN_5845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5847 = 7'h2d == _myNewVec_83_T_3[6:0] ? myVec_45 : _GEN_5846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5848 = 7'h2e == _myNewVec_83_T_3[6:0] ? myVec_46 : _GEN_5847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5849 = 7'h2f == _myNewVec_83_T_3[6:0] ? myVec_47 : _GEN_5848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5850 = 7'h30 == _myNewVec_83_T_3[6:0] ? myVec_48 : _GEN_5849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5851 = 7'h31 == _myNewVec_83_T_3[6:0] ? myVec_49 : _GEN_5850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5852 = 7'h32 == _myNewVec_83_T_3[6:0] ? myVec_50 : _GEN_5851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5853 = 7'h33 == _myNewVec_83_T_3[6:0] ? myVec_51 : _GEN_5852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5854 = 7'h34 == _myNewVec_83_T_3[6:0] ? myVec_52 : _GEN_5853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5855 = 7'h35 == _myNewVec_83_T_3[6:0] ? myVec_53 : _GEN_5854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5856 = 7'h36 == _myNewVec_83_T_3[6:0] ? myVec_54 : _GEN_5855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5857 = 7'h37 == _myNewVec_83_T_3[6:0] ? myVec_55 : _GEN_5856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5858 = 7'h38 == _myNewVec_83_T_3[6:0] ? myVec_56 : _GEN_5857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5859 = 7'h39 == _myNewVec_83_T_3[6:0] ? myVec_57 : _GEN_5858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5860 = 7'h3a == _myNewVec_83_T_3[6:0] ? myVec_58 : _GEN_5859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5861 = 7'h3b == _myNewVec_83_T_3[6:0] ? myVec_59 : _GEN_5860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5862 = 7'h3c == _myNewVec_83_T_3[6:0] ? myVec_60 : _GEN_5861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5863 = 7'h3d == _myNewVec_83_T_3[6:0] ? myVec_61 : _GEN_5862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5864 = 7'h3e == _myNewVec_83_T_3[6:0] ? myVec_62 : _GEN_5863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5865 = 7'h3f == _myNewVec_83_T_3[6:0] ? myVec_63 : _GEN_5864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5866 = 7'h40 == _myNewVec_83_T_3[6:0] ? myVec_64 : _GEN_5865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5867 = 7'h41 == _myNewVec_83_T_3[6:0] ? myVec_65 : _GEN_5866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5868 = 7'h42 == _myNewVec_83_T_3[6:0] ? myVec_66 : _GEN_5867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5869 = 7'h43 == _myNewVec_83_T_3[6:0] ? myVec_67 : _GEN_5868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5870 = 7'h44 == _myNewVec_83_T_3[6:0] ? myVec_68 : _GEN_5869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5871 = 7'h45 == _myNewVec_83_T_3[6:0] ? myVec_69 : _GEN_5870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5872 = 7'h46 == _myNewVec_83_T_3[6:0] ? myVec_70 : _GEN_5871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5873 = 7'h47 == _myNewVec_83_T_3[6:0] ? myVec_71 : _GEN_5872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5874 = 7'h48 == _myNewVec_83_T_3[6:0] ? myVec_72 : _GEN_5873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5875 = 7'h49 == _myNewVec_83_T_3[6:0] ? myVec_73 : _GEN_5874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5876 = 7'h4a == _myNewVec_83_T_3[6:0] ? myVec_74 : _GEN_5875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5877 = 7'h4b == _myNewVec_83_T_3[6:0] ? myVec_75 : _GEN_5876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5878 = 7'h4c == _myNewVec_83_T_3[6:0] ? myVec_76 : _GEN_5877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5879 = 7'h4d == _myNewVec_83_T_3[6:0] ? myVec_77 : _GEN_5878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5880 = 7'h4e == _myNewVec_83_T_3[6:0] ? myVec_78 : _GEN_5879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5881 = 7'h4f == _myNewVec_83_T_3[6:0] ? myVec_79 : _GEN_5880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5882 = 7'h50 == _myNewVec_83_T_3[6:0] ? myVec_80 : _GEN_5881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5883 = 7'h51 == _myNewVec_83_T_3[6:0] ? myVec_81 : _GEN_5882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5884 = 7'h52 == _myNewVec_83_T_3[6:0] ? myVec_82 : _GEN_5883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5885 = 7'h53 == _myNewVec_83_T_3[6:0] ? myVec_83 : _GEN_5884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5886 = 7'h54 == _myNewVec_83_T_3[6:0] ? myVec_84 : _GEN_5885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5887 = 7'h55 == _myNewVec_83_T_3[6:0] ? myVec_85 : _GEN_5886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5888 = 7'h56 == _myNewVec_83_T_3[6:0] ? myVec_86 : _GEN_5887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5889 = 7'h57 == _myNewVec_83_T_3[6:0] ? myVec_87 : _GEN_5888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5890 = 7'h58 == _myNewVec_83_T_3[6:0] ? myVec_88 : _GEN_5889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5891 = 7'h59 == _myNewVec_83_T_3[6:0] ? myVec_89 : _GEN_5890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5892 = 7'h5a == _myNewVec_83_T_3[6:0] ? myVec_90 : _GEN_5891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5893 = 7'h5b == _myNewVec_83_T_3[6:0] ? myVec_91 : _GEN_5892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5894 = 7'h5c == _myNewVec_83_T_3[6:0] ? myVec_92 : _GEN_5893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5895 = 7'h5d == _myNewVec_83_T_3[6:0] ? myVec_93 : _GEN_5894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5896 = 7'h5e == _myNewVec_83_T_3[6:0] ? myVec_94 : _GEN_5895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5897 = 7'h5f == _myNewVec_83_T_3[6:0] ? myVec_95 : _GEN_5896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5898 = 7'h60 == _myNewVec_83_T_3[6:0] ? myVec_96 : _GEN_5897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5899 = 7'h61 == _myNewVec_83_T_3[6:0] ? myVec_97 : _GEN_5898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5900 = 7'h62 == _myNewVec_83_T_3[6:0] ? myVec_98 : _GEN_5899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5901 = 7'h63 == _myNewVec_83_T_3[6:0] ? myVec_99 : _GEN_5900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5902 = 7'h64 == _myNewVec_83_T_3[6:0] ? myVec_100 : _GEN_5901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5903 = 7'h65 == _myNewVec_83_T_3[6:0] ? myVec_101 : _GEN_5902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5904 = 7'h66 == _myNewVec_83_T_3[6:0] ? myVec_102 : _GEN_5903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5905 = 7'h67 == _myNewVec_83_T_3[6:0] ? myVec_103 : _GEN_5904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5906 = 7'h68 == _myNewVec_83_T_3[6:0] ? myVec_104 : _GEN_5905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5907 = 7'h69 == _myNewVec_83_T_3[6:0] ? myVec_105 : _GEN_5906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5908 = 7'h6a == _myNewVec_83_T_3[6:0] ? myVec_106 : _GEN_5907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5909 = 7'h6b == _myNewVec_83_T_3[6:0] ? myVec_107 : _GEN_5908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5910 = 7'h6c == _myNewVec_83_T_3[6:0] ? myVec_108 : _GEN_5909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5911 = 7'h6d == _myNewVec_83_T_3[6:0] ? myVec_109 : _GEN_5910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5912 = 7'h6e == _myNewVec_83_T_3[6:0] ? myVec_110 : _GEN_5911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5913 = 7'h6f == _myNewVec_83_T_3[6:0] ? myVec_111 : _GEN_5912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5914 = 7'h70 == _myNewVec_83_T_3[6:0] ? myVec_112 : _GEN_5913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5915 = 7'h71 == _myNewVec_83_T_3[6:0] ? myVec_113 : _GEN_5914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5916 = 7'h72 == _myNewVec_83_T_3[6:0] ? myVec_114 : _GEN_5915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5917 = 7'h73 == _myNewVec_83_T_3[6:0] ? myVec_115 : _GEN_5916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5918 = 7'h74 == _myNewVec_83_T_3[6:0] ? myVec_116 : _GEN_5917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5919 = 7'h75 == _myNewVec_83_T_3[6:0] ? myVec_117 : _GEN_5918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5920 = 7'h76 == _myNewVec_83_T_3[6:0] ? myVec_118 : _GEN_5919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5921 = 7'h77 == _myNewVec_83_T_3[6:0] ? myVec_119 : _GEN_5920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5922 = 7'h78 == _myNewVec_83_T_3[6:0] ? myVec_120 : _GEN_5921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5923 = 7'h79 == _myNewVec_83_T_3[6:0] ? myVec_121 : _GEN_5922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5924 = 7'h7a == _myNewVec_83_T_3[6:0] ? myVec_122 : _GEN_5923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5925 = 7'h7b == _myNewVec_83_T_3[6:0] ? myVec_123 : _GEN_5924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5926 = 7'h7c == _myNewVec_83_T_3[6:0] ? myVec_124 : _GEN_5925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5927 = 7'h7d == _myNewVec_83_T_3[6:0] ? myVec_125 : _GEN_5926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5928 = 7'h7e == _myNewVec_83_T_3[6:0] ? myVec_126 : _GEN_5927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_83 = 7'h7f == _myNewVec_83_T_3[6:0] ? myVec_127 : _GEN_5928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_82_T_3 = _myNewVec_127_T_1 + 16'h2d; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_5931 = 7'h1 == _myNewVec_82_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5932 = 7'h2 == _myNewVec_82_T_3[6:0] ? myVec_2 : _GEN_5931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5933 = 7'h3 == _myNewVec_82_T_3[6:0] ? myVec_3 : _GEN_5932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5934 = 7'h4 == _myNewVec_82_T_3[6:0] ? myVec_4 : _GEN_5933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5935 = 7'h5 == _myNewVec_82_T_3[6:0] ? myVec_5 : _GEN_5934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5936 = 7'h6 == _myNewVec_82_T_3[6:0] ? myVec_6 : _GEN_5935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5937 = 7'h7 == _myNewVec_82_T_3[6:0] ? myVec_7 : _GEN_5936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5938 = 7'h8 == _myNewVec_82_T_3[6:0] ? myVec_8 : _GEN_5937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5939 = 7'h9 == _myNewVec_82_T_3[6:0] ? myVec_9 : _GEN_5938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5940 = 7'ha == _myNewVec_82_T_3[6:0] ? myVec_10 : _GEN_5939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5941 = 7'hb == _myNewVec_82_T_3[6:0] ? myVec_11 : _GEN_5940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5942 = 7'hc == _myNewVec_82_T_3[6:0] ? myVec_12 : _GEN_5941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5943 = 7'hd == _myNewVec_82_T_3[6:0] ? myVec_13 : _GEN_5942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5944 = 7'he == _myNewVec_82_T_3[6:0] ? myVec_14 : _GEN_5943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5945 = 7'hf == _myNewVec_82_T_3[6:0] ? myVec_15 : _GEN_5944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5946 = 7'h10 == _myNewVec_82_T_3[6:0] ? myVec_16 : _GEN_5945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5947 = 7'h11 == _myNewVec_82_T_3[6:0] ? myVec_17 : _GEN_5946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5948 = 7'h12 == _myNewVec_82_T_3[6:0] ? myVec_18 : _GEN_5947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5949 = 7'h13 == _myNewVec_82_T_3[6:0] ? myVec_19 : _GEN_5948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5950 = 7'h14 == _myNewVec_82_T_3[6:0] ? myVec_20 : _GEN_5949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5951 = 7'h15 == _myNewVec_82_T_3[6:0] ? myVec_21 : _GEN_5950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5952 = 7'h16 == _myNewVec_82_T_3[6:0] ? myVec_22 : _GEN_5951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5953 = 7'h17 == _myNewVec_82_T_3[6:0] ? myVec_23 : _GEN_5952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5954 = 7'h18 == _myNewVec_82_T_3[6:0] ? myVec_24 : _GEN_5953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5955 = 7'h19 == _myNewVec_82_T_3[6:0] ? myVec_25 : _GEN_5954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5956 = 7'h1a == _myNewVec_82_T_3[6:0] ? myVec_26 : _GEN_5955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5957 = 7'h1b == _myNewVec_82_T_3[6:0] ? myVec_27 : _GEN_5956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5958 = 7'h1c == _myNewVec_82_T_3[6:0] ? myVec_28 : _GEN_5957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5959 = 7'h1d == _myNewVec_82_T_3[6:0] ? myVec_29 : _GEN_5958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5960 = 7'h1e == _myNewVec_82_T_3[6:0] ? myVec_30 : _GEN_5959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5961 = 7'h1f == _myNewVec_82_T_3[6:0] ? myVec_31 : _GEN_5960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5962 = 7'h20 == _myNewVec_82_T_3[6:0] ? myVec_32 : _GEN_5961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5963 = 7'h21 == _myNewVec_82_T_3[6:0] ? myVec_33 : _GEN_5962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5964 = 7'h22 == _myNewVec_82_T_3[6:0] ? myVec_34 : _GEN_5963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5965 = 7'h23 == _myNewVec_82_T_3[6:0] ? myVec_35 : _GEN_5964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5966 = 7'h24 == _myNewVec_82_T_3[6:0] ? myVec_36 : _GEN_5965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5967 = 7'h25 == _myNewVec_82_T_3[6:0] ? myVec_37 : _GEN_5966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5968 = 7'h26 == _myNewVec_82_T_3[6:0] ? myVec_38 : _GEN_5967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5969 = 7'h27 == _myNewVec_82_T_3[6:0] ? myVec_39 : _GEN_5968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5970 = 7'h28 == _myNewVec_82_T_3[6:0] ? myVec_40 : _GEN_5969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5971 = 7'h29 == _myNewVec_82_T_3[6:0] ? myVec_41 : _GEN_5970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5972 = 7'h2a == _myNewVec_82_T_3[6:0] ? myVec_42 : _GEN_5971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5973 = 7'h2b == _myNewVec_82_T_3[6:0] ? myVec_43 : _GEN_5972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5974 = 7'h2c == _myNewVec_82_T_3[6:0] ? myVec_44 : _GEN_5973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5975 = 7'h2d == _myNewVec_82_T_3[6:0] ? myVec_45 : _GEN_5974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5976 = 7'h2e == _myNewVec_82_T_3[6:0] ? myVec_46 : _GEN_5975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5977 = 7'h2f == _myNewVec_82_T_3[6:0] ? myVec_47 : _GEN_5976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5978 = 7'h30 == _myNewVec_82_T_3[6:0] ? myVec_48 : _GEN_5977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5979 = 7'h31 == _myNewVec_82_T_3[6:0] ? myVec_49 : _GEN_5978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5980 = 7'h32 == _myNewVec_82_T_3[6:0] ? myVec_50 : _GEN_5979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5981 = 7'h33 == _myNewVec_82_T_3[6:0] ? myVec_51 : _GEN_5980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5982 = 7'h34 == _myNewVec_82_T_3[6:0] ? myVec_52 : _GEN_5981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5983 = 7'h35 == _myNewVec_82_T_3[6:0] ? myVec_53 : _GEN_5982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5984 = 7'h36 == _myNewVec_82_T_3[6:0] ? myVec_54 : _GEN_5983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5985 = 7'h37 == _myNewVec_82_T_3[6:0] ? myVec_55 : _GEN_5984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5986 = 7'h38 == _myNewVec_82_T_3[6:0] ? myVec_56 : _GEN_5985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5987 = 7'h39 == _myNewVec_82_T_3[6:0] ? myVec_57 : _GEN_5986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5988 = 7'h3a == _myNewVec_82_T_3[6:0] ? myVec_58 : _GEN_5987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5989 = 7'h3b == _myNewVec_82_T_3[6:0] ? myVec_59 : _GEN_5988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5990 = 7'h3c == _myNewVec_82_T_3[6:0] ? myVec_60 : _GEN_5989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5991 = 7'h3d == _myNewVec_82_T_3[6:0] ? myVec_61 : _GEN_5990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5992 = 7'h3e == _myNewVec_82_T_3[6:0] ? myVec_62 : _GEN_5991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5993 = 7'h3f == _myNewVec_82_T_3[6:0] ? myVec_63 : _GEN_5992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5994 = 7'h40 == _myNewVec_82_T_3[6:0] ? myVec_64 : _GEN_5993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5995 = 7'h41 == _myNewVec_82_T_3[6:0] ? myVec_65 : _GEN_5994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5996 = 7'h42 == _myNewVec_82_T_3[6:0] ? myVec_66 : _GEN_5995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5997 = 7'h43 == _myNewVec_82_T_3[6:0] ? myVec_67 : _GEN_5996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5998 = 7'h44 == _myNewVec_82_T_3[6:0] ? myVec_68 : _GEN_5997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_5999 = 7'h45 == _myNewVec_82_T_3[6:0] ? myVec_69 : _GEN_5998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6000 = 7'h46 == _myNewVec_82_T_3[6:0] ? myVec_70 : _GEN_5999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6001 = 7'h47 == _myNewVec_82_T_3[6:0] ? myVec_71 : _GEN_6000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6002 = 7'h48 == _myNewVec_82_T_3[6:0] ? myVec_72 : _GEN_6001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6003 = 7'h49 == _myNewVec_82_T_3[6:0] ? myVec_73 : _GEN_6002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6004 = 7'h4a == _myNewVec_82_T_3[6:0] ? myVec_74 : _GEN_6003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6005 = 7'h4b == _myNewVec_82_T_3[6:0] ? myVec_75 : _GEN_6004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6006 = 7'h4c == _myNewVec_82_T_3[6:0] ? myVec_76 : _GEN_6005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6007 = 7'h4d == _myNewVec_82_T_3[6:0] ? myVec_77 : _GEN_6006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6008 = 7'h4e == _myNewVec_82_T_3[6:0] ? myVec_78 : _GEN_6007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6009 = 7'h4f == _myNewVec_82_T_3[6:0] ? myVec_79 : _GEN_6008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6010 = 7'h50 == _myNewVec_82_T_3[6:0] ? myVec_80 : _GEN_6009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6011 = 7'h51 == _myNewVec_82_T_3[6:0] ? myVec_81 : _GEN_6010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6012 = 7'h52 == _myNewVec_82_T_3[6:0] ? myVec_82 : _GEN_6011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6013 = 7'h53 == _myNewVec_82_T_3[6:0] ? myVec_83 : _GEN_6012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6014 = 7'h54 == _myNewVec_82_T_3[6:0] ? myVec_84 : _GEN_6013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6015 = 7'h55 == _myNewVec_82_T_3[6:0] ? myVec_85 : _GEN_6014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6016 = 7'h56 == _myNewVec_82_T_3[6:0] ? myVec_86 : _GEN_6015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6017 = 7'h57 == _myNewVec_82_T_3[6:0] ? myVec_87 : _GEN_6016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6018 = 7'h58 == _myNewVec_82_T_3[6:0] ? myVec_88 : _GEN_6017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6019 = 7'h59 == _myNewVec_82_T_3[6:0] ? myVec_89 : _GEN_6018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6020 = 7'h5a == _myNewVec_82_T_3[6:0] ? myVec_90 : _GEN_6019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6021 = 7'h5b == _myNewVec_82_T_3[6:0] ? myVec_91 : _GEN_6020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6022 = 7'h5c == _myNewVec_82_T_3[6:0] ? myVec_92 : _GEN_6021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6023 = 7'h5d == _myNewVec_82_T_3[6:0] ? myVec_93 : _GEN_6022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6024 = 7'h5e == _myNewVec_82_T_3[6:0] ? myVec_94 : _GEN_6023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6025 = 7'h5f == _myNewVec_82_T_3[6:0] ? myVec_95 : _GEN_6024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6026 = 7'h60 == _myNewVec_82_T_3[6:0] ? myVec_96 : _GEN_6025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6027 = 7'h61 == _myNewVec_82_T_3[6:0] ? myVec_97 : _GEN_6026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6028 = 7'h62 == _myNewVec_82_T_3[6:0] ? myVec_98 : _GEN_6027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6029 = 7'h63 == _myNewVec_82_T_3[6:0] ? myVec_99 : _GEN_6028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6030 = 7'h64 == _myNewVec_82_T_3[6:0] ? myVec_100 : _GEN_6029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6031 = 7'h65 == _myNewVec_82_T_3[6:0] ? myVec_101 : _GEN_6030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6032 = 7'h66 == _myNewVec_82_T_3[6:0] ? myVec_102 : _GEN_6031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6033 = 7'h67 == _myNewVec_82_T_3[6:0] ? myVec_103 : _GEN_6032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6034 = 7'h68 == _myNewVec_82_T_3[6:0] ? myVec_104 : _GEN_6033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6035 = 7'h69 == _myNewVec_82_T_3[6:0] ? myVec_105 : _GEN_6034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6036 = 7'h6a == _myNewVec_82_T_3[6:0] ? myVec_106 : _GEN_6035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6037 = 7'h6b == _myNewVec_82_T_3[6:0] ? myVec_107 : _GEN_6036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6038 = 7'h6c == _myNewVec_82_T_3[6:0] ? myVec_108 : _GEN_6037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6039 = 7'h6d == _myNewVec_82_T_3[6:0] ? myVec_109 : _GEN_6038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6040 = 7'h6e == _myNewVec_82_T_3[6:0] ? myVec_110 : _GEN_6039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6041 = 7'h6f == _myNewVec_82_T_3[6:0] ? myVec_111 : _GEN_6040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6042 = 7'h70 == _myNewVec_82_T_3[6:0] ? myVec_112 : _GEN_6041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6043 = 7'h71 == _myNewVec_82_T_3[6:0] ? myVec_113 : _GEN_6042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6044 = 7'h72 == _myNewVec_82_T_3[6:0] ? myVec_114 : _GEN_6043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6045 = 7'h73 == _myNewVec_82_T_3[6:0] ? myVec_115 : _GEN_6044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6046 = 7'h74 == _myNewVec_82_T_3[6:0] ? myVec_116 : _GEN_6045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6047 = 7'h75 == _myNewVec_82_T_3[6:0] ? myVec_117 : _GEN_6046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6048 = 7'h76 == _myNewVec_82_T_3[6:0] ? myVec_118 : _GEN_6047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6049 = 7'h77 == _myNewVec_82_T_3[6:0] ? myVec_119 : _GEN_6048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6050 = 7'h78 == _myNewVec_82_T_3[6:0] ? myVec_120 : _GEN_6049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6051 = 7'h79 == _myNewVec_82_T_3[6:0] ? myVec_121 : _GEN_6050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6052 = 7'h7a == _myNewVec_82_T_3[6:0] ? myVec_122 : _GEN_6051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6053 = 7'h7b == _myNewVec_82_T_3[6:0] ? myVec_123 : _GEN_6052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6054 = 7'h7c == _myNewVec_82_T_3[6:0] ? myVec_124 : _GEN_6053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6055 = 7'h7d == _myNewVec_82_T_3[6:0] ? myVec_125 : _GEN_6054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6056 = 7'h7e == _myNewVec_82_T_3[6:0] ? myVec_126 : _GEN_6055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_82 = 7'h7f == _myNewVec_82_T_3[6:0] ? myVec_127 : _GEN_6056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_81_T_3 = _myNewVec_127_T_1 + 16'h2e; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_6059 = 7'h1 == _myNewVec_81_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6060 = 7'h2 == _myNewVec_81_T_3[6:0] ? myVec_2 : _GEN_6059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6061 = 7'h3 == _myNewVec_81_T_3[6:0] ? myVec_3 : _GEN_6060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6062 = 7'h4 == _myNewVec_81_T_3[6:0] ? myVec_4 : _GEN_6061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6063 = 7'h5 == _myNewVec_81_T_3[6:0] ? myVec_5 : _GEN_6062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6064 = 7'h6 == _myNewVec_81_T_3[6:0] ? myVec_6 : _GEN_6063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6065 = 7'h7 == _myNewVec_81_T_3[6:0] ? myVec_7 : _GEN_6064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6066 = 7'h8 == _myNewVec_81_T_3[6:0] ? myVec_8 : _GEN_6065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6067 = 7'h9 == _myNewVec_81_T_3[6:0] ? myVec_9 : _GEN_6066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6068 = 7'ha == _myNewVec_81_T_3[6:0] ? myVec_10 : _GEN_6067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6069 = 7'hb == _myNewVec_81_T_3[6:0] ? myVec_11 : _GEN_6068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6070 = 7'hc == _myNewVec_81_T_3[6:0] ? myVec_12 : _GEN_6069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6071 = 7'hd == _myNewVec_81_T_3[6:0] ? myVec_13 : _GEN_6070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6072 = 7'he == _myNewVec_81_T_3[6:0] ? myVec_14 : _GEN_6071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6073 = 7'hf == _myNewVec_81_T_3[6:0] ? myVec_15 : _GEN_6072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6074 = 7'h10 == _myNewVec_81_T_3[6:0] ? myVec_16 : _GEN_6073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6075 = 7'h11 == _myNewVec_81_T_3[6:0] ? myVec_17 : _GEN_6074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6076 = 7'h12 == _myNewVec_81_T_3[6:0] ? myVec_18 : _GEN_6075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6077 = 7'h13 == _myNewVec_81_T_3[6:0] ? myVec_19 : _GEN_6076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6078 = 7'h14 == _myNewVec_81_T_3[6:0] ? myVec_20 : _GEN_6077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6079 = 7'h15 == _myNewVec_81_T_3[6:0] ? myVec_21 : _GEN_6078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6080 = 7'h16 == _myNewVec_81_T_3[6:0] ? myVec_22 : _GEN_6079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6081 = 7'h17 == _myNewVec_81_T_3[6:0] ? myVec_23 : _GEN_6080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6082 = 7'h18 == _myNewVec_81_T_3[6:0] ? myVec_24 : _GEN_6081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6083 = 7'h19 == _myNewVec_81_T_3[6:0] ? myVec_25 : _GEN_6082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6084 = 7'h1a == _myNewVec_81_T_3[6:0] ? myVec_26 : _GEN_6083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6085 = 7'h1b == _myNewVec_81_T_3[6:0] ? myVec_27 : _GEN_6084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6086 = 7'h1c == _myNewVec_81_T_3[6:0] ? myVec_28 : _GEN_6085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6087 = 7'h1d == _myNewVec_81_T_3[6:0] ? myVec_29 : _GEN_6086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6088 = 7'h1e == _myNewVec_81_T_3[6:0] ? myVec_30 : _GEN_6087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6089 = 7'h1f == _myNewVec_81_T_3[6:0] ? myVec_31 : _GEN_6088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6090 = 7'h20 == _myNewVec_81_T_3[6:0] ? myVec_32 : _GEN_6089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6091 = 7'h21 == _myNewVec_81_T_3[6:0] ? myVec_33 : _GEN_6090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6092 = 7'h22 == _myNewVec_81_T_3[6:0] ? myVec_34 : _GEN_6091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6093 = 7'h23 == _myNewVec_81_T_3[6:0] ? myVec_35 : _GEN_6092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6094 = 7'h24 == _myNewVec_81_T_3[6:0] ? myVec_36 : _GEN_6093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6095 = 7'h25 == _myNewVec_81_T_3[6:0] ? myVec_37 : _GEN_6094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6096 = 7'h26 == _myNewVec_81_T_3[6:0] ? myVec_38 : _GEN_6095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6097 = 7'h27 == _myNewVec_81_T_3[6:0] ? myVec_39 : _GEN_6096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6098 = 7'h28 == _myNewVec_81_T_3[6:0] ? myVec_40 : _GEN_6097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6099 = 7'h29 == _myNewVec_81_T_3[6:0] ? myVec_41 : _GEN_6098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6100 = 7'h2a == _myNewVec_81_T_3[6:0] ? myVec_42 : _GEN_6099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6101 = 7'h2b == _myNewVec_81_T_3[6:0] ? myVec_43 : _GEN_6100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6102 = 7'h2c == _myNewVec_81_T_3[6:0] ? myVec_44 : _GEN_6101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6103 = 7'h2d == _myNewVec_81_T_3[6:0] ? myVec_45 : _GEN_6102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6104 = 7'h2e == _myNewVec_81_T_3[6:0] ? myVec_46 : _GEN_6103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6105 = 7'h2f == _myNewVec_81_T_3[6:0] ? myVec_47 : _GEN_6104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6106 = 7'h30 == _myNewVec_81_T_3[6:0] ? myVec_48 : _GEN_6105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6107 = 7'h31 == _myNewVec_81_T_3[6:0] ? myVec_49 : _GEN_6106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6108 = 7'h32 == _myNewVec_81_T_3[6:0] ? myVec_50 : _GEN_6107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6109 = 7'h33 == _myNewVec_81_T_3[6:0] ? myVec_51 : _GEN_6108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6110 = 7'h34 == _myNewVec_81_T_3[6:0] ? myVec_52 : _GEN_6109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6111 = 7'h35 == _myNewVec_81_T_3[6:0] ? myVec_53 : _GEN_6110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6112 = 7'h36 == _myNewVec_81_T_3[6:0] ? myVec_54 : _GEN_6111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6113 = 7'h37 == _myNewVec_81_T_3[6:0] ? myVec_55 : _GEN_6112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6114 = 7'h38 == _myNewVec_81_T_3[6:0] ? myVec_56 : _GEN_6113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6115 = 7'h39 == _myNewVec_81_T_3[6:0] ? myVec_57 : _GEN_6114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6116 = 7'h3a == _myNewVec_81_T_3[6:0] ? myVec_58 : _GEN_6115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6117 = 7'h3b == _myNewVec_81_T_3[6:0] ? myVec_59 : _GEN_6116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6118 = 7'h3c == _myNewVec_81_T_3[6:0] ? myVec_60 : _GEN_6117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6119 = 7'h3d == _myNewVec_81_T_3[6:0] ? myVec_61 : _GEN_6118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6120 = 7'h3e == _myNewVec_81_T_3[6:0] ? myVec_62 : _GEN_6119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6121 = 7'h3f == _myNewVec_81_T_3[6:0] ? myVec_63 : _GEN_6120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6122 = 7'h40 == _myNewVec_81_T_3[6:0] ? myVec_64 : _GEN_6121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6123 = 7'h41 == _myNewVec_81_T_3[6:0] ? myVec_65 : _GEN_6122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6124 = 7'h42 == _myNewVec_81_T_3[6:0] ? myVec_66 : _GEN_6123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6125 = 7'h43 == _myNewVec_81_T_3[6:0] ? myVec_67 : _GEN_6124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6126 = 7'h44 == _myNewVec_81_T_3[6:0] ? myVec_68 : _GEN_6125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6127 = 7'h45 == _myNewVec_81_T_3[6:0] ? myVec_69 : _GEN_6126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6128 = 7'h46 == _myNewVec_81_T_3[6:0] ? myVec_70 : _GEN_6127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6129 = 7'h47 == _myNewVec_81_T_3[6:0] ? myVec_71 : _GEN_6128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6130 = 7'h48 == _myNewVec_81_T_3[6:0] ? myVec_72 : _GEN_6129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6131 = 7'h49 == _myNewVec_81_T_3[6:0] ? myVec_73 : _GEN_6130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6132 = 7'h4a == _myNewVec_81_T_3[6:0] ? myVec_74 : _GEN_6131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6133 = 7'h4b == _myNewVec_81_T_3[6:0] ? myVec_75 : _GEN_6132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6134 = 7'h4c == _myNewVec_81_T_3[6:0] ? myVec_76 : _GEN_6133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6135 = 7'h4d == _myNewVec_81_T_3[6:0] ? myVec_77 : _GEN_6134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6136 = 7'h4e == _myNewVec_81_T_3[6:0] ? myVec_78 : _GEN_6135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6137 = 7'h4f == _myNewVec_81_T_3[6:0] ? myVec_79 : _GEN_6136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6138 = 7'h50 == _myNewVec_81_T_3[6:0] ? myVec_80 : _GEN_6137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6139 = 7'h51 == _myNewVec_81_T_3[6:0] ? myVec_81 : _GEN_6138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6140 = 7'h52 == _myNewVec_81_T_3[6:0] ? myVec_82 : _GEN_6139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6141 = 7'h53 == _myNewVec_81_T_3[6:0] ? myVec_83 : _GEN_6140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6142 = 7'h54 == _myNewVec_81_T_3[6:0] ? myVec_84 : _GEN_6141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6143 = 7'h55 == _myNewVec_81_T_3[6:0] ? myVec_85 : _GEN_6142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6144 = 7'h56 == _myNewVec_81_T_3[6:0] ? myVec_86 : _GEN_6143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6145 = 7'h57 == _myNewVec_81_T_3[6:0] ? myVec_87 : _GEN_6144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6146 = 7'h58 == _myNewVec_81_T_3[6:0] ? myVec_88 : _GEN_6145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6147 = 7'h59 == _myNewVec_81_T_3[6:0] ? myVec_89 : _GEN_6146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6148 = 7'h5a == _myNewVec_81_T_3[6:0] ? myVec_90 : _GEN_6147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6149 = 7'h5b == _myNewVec_81_T_3[6:0] ? myVec_91 : _GEN_6148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6150 = 7'h5c == _myNewVec_81_T_3[6:0] ? myVec_92 : _GEN_6149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6151 = 7'h5d == _myNewVec_81_T_3[6:0] ? myVec_93 : _GEN_6150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6152 = 7'h5e == _myNewVec_81_T_3[6:0] ? myVec_94 : _GEN_6151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6153 = 7'h5f == _myNewVec_81_T_3[6:0] ? myVec_95 : _GEN_6152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6154 = 7'h60 == _myNewVec_81_T_3[6:0] ? myVec_96 : _GEN_6153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6155 = 7'h61 == _myNewVec_81_T_3[6:0] ? myVec_97 : _GEN_6154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6156 = 7'h62 == _myNewVec_81_T_3[6:0] ? myVec_98 : _GEN_6155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6157 = 7'h63 == _myNewVec_81_T_3[6:0] ? myVec_99 : _GEN_6156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6158 = 7'h64 == _myNewVec_81_T_3[6:0] ? myVec_100 : _GEN_6157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6159 = 7'h65 == _myNewVec_81_T_3[6:0] ? myVec_101 : _GEN_6158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6160 = 7'h66 == _myNewVec_81_T_3[6:0] ? myVec_102 : _GEN_6159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6161 = 7'h67 == _myNewVec_81_T_3[6:0] ? myVec_103 : _GEN_6160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6162 = 7'h68 == _myNewVec_81_T_3[6:0] ? myVec_104 : _GEN_6161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6163 = 7'h69 == _myNewVec_81_T_3[6:0] ? myVec_105 : _GEN_6162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6164 = 7'h6a == _myNewVec_81_T_3[6:0] ? myVec_106 : _GEN_6163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6165 = 7'h6b == _myNewVec_81_T_3[6:0] ? myVec_107 : _GEN_6164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6166 = 7'h6c == _myNewVec_81_T_3[6:0] ? myVec_108 : _GEN_6165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6167 = 7'h6d == _myNewVec_81_T_3[6:0] ? myVec_109 : _GEN_6166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6168 = 7'h6e == _myNewVec_81_T_3[6:0] ? myVec_110 : _GEN_6167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6169 = 7'h6f == _myNewVec_81_T_3[6:0] ? myVec_111 : _GEN_6168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6170 = 7'h70 == _myNewVec_81_T_3[6:0] ? myVec_112 : _GEN_6169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6171 = 7'h71 == _myNewVec_81_T_3[6:0] ? myVec_113 : _GEN_6170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6172 = 7'h72 == _myNewVec_81_T_3[6:0] ? myVec_114 : _GEN_6171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6173 = 7'h73 == _myNewVec_81_T_3[6:0] ? myVec_115 : _GEN_6172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6174 = 7'h74 == _myNewVec_81_T_3[6:0] ? myVec_116 : _GEN_6173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6175 = 7'h75 == _myNewVec_81_T_3[6:0] ? myVec_117 : _GEN_6174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6176 = 7'h76 == _myNewVec_81_T_3[6:0] ? myVec_118 : _GEN_6175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6177 = 7'h77 == _myNewVec_81_T_3[6:0] ? myVec_119 : _GEN_6176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6178 = 7'h78 == _myNewVec_81_T_3[6:0] ? myVec_120 : _GEN_6177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6179 = 7'h79 == _myNewVec_81_T_3[6:0] ? myVec_121 : _GEN_6178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6180 = 7'h7a == _myNewVec_81_T_3[6:0] ? myVec_122 : _GEN_6179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6181 = 7'h7b == _myNewVec_81_T_3[6:0] ? myVec_123 : _GEN_6180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6182 = 7'h7c == _myNewVec_81_T_3[6:0] ? myVec_124 : _GEN_6181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6183 = 7'h7d == _myNewVec_81_T_3[6:0] ? myVec_125 : _GEN_6182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6184 = 7'h7e == _myNewVec_81_T_3[6:0] ? myVec_126 : _GEN_6183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_81 = 7'h7f == _myNewVec_81_T_3[6:0] ? myVec_127 : _GEN_6184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_80_T_3 = _myNewVec_127_T_1 + 16'h2f; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_6187 = 7'h1 == _myNewVec_80_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6188 = 7'h2 == _myNewVec_80_T_3[6:0] ? myVec_2 : _GEN_6187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6189 = 7'h3 == _myNewVec_80_T_3[6:0] ? myVec_3 : _GEN_6188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6190 = 7'h4 == _myNewVec_80_T_3[6:0] ? myVec_4 : _GEN_6189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6191 = 7'h5 == _myNewVec_80_T_3[6:0] ? myVec_5 : _GEN_6190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6192 = 7'h6 == _myNewVec_80_T_3[6:0] ? myVec_6 : _GEN_6191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6193 = 7'h7 == _myNewVec_80_T_3[6:0] ? myVec_7 : _GEN_6192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6194 = 7'h8 == _myNewVec_80_T_3[6:0] ? myVec_8 : _GEN_6193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6195 = 7'h9 == _myNewVec_80_T_3[6:0] ? myVec_9 : _GEN_6194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6196 = 7'ha == _myNewVec_80_T_3[6:0] ? myVec_10 : _GEN_6195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6197 = 7'hb == _myNewVec_80_T_3[6:0] ? myVec_11 : _GEN_6196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6198 = 7'hc == _myNewVec_80_T_3[6:0] ? myVec_12 : _GEN_6197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6199 = 7'hd == _myNewVec_80_T_3[6:0] ? myVec_13 : _GEN_6198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6200 = 7'he == _myNewVec_80_T_3[6:0] ? myVec_14 : _GEN_6199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6201 = 7'hf == _myNewVec_80_T_3[6:0] ? myVec_15 : _GEN_6200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6202 = 7'h10 == _myNewVec_80_T_3[6:0] ? myVec_16 : _GEN_6201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6203 = 7'h11 == _myNewVec_80_T_3[6:0] ? myVec_17 : _GEN_6202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6204 = 7'h12 == _myNewVec_80_T_3[6:0] ? myVec_18 : _GEN_6203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6205 = 7'h13 == _myNewVec_80_T_3[6:0] ? myVec_19 : _GEN_6204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6206 = 7'h14 == _myNewVec_80_T_3[6:0] ? myVec_20 : _GEN_6205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6207 = 7'h15 == _myNewVec_80_T_3[6:0] ? myVec_21 : _GEN_6206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6208 = 7'h16 == _myNewVec_80_T_3[6:0] ? myVec_22 : _GEN_6207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6209 = 7'h17 == _myNewVec_80_T_3[6:0] ? myVec_23 : _GEN_6208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6210 = 7'h18 == _myNewVec_80_T_3[6:0] ? myVec_24 : _GEN_6209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6211 = 7'h19 == _myNewVec_80_T_3[6:0] ? myVec_25 : _GEN_6210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6212 = 7'h1a == _myNewVec_80_T_3[6:0] ? myVec_26 : _GEN_6211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6213 = 7'h1b == _myNewVec_80_T_3[6:0] ? myVec_27 : _GEN_6212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6214 = 7'h1c == _myNewVec_80_T_3[6:0] ? myVec_28 : _GEN_6213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6215 = 7'h1d == _myNewVec_80_T_3[6:0] ? myVec_29 : _GEN_6214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6216 = 7'h1e == _myNewVec_80_T_3[6:0] ? myVec_30 : _GEN_6215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6217 = 7'h1f == _myNewVec_80_T_3[6:0] ? myVec_31 : _GEN_6216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6218 = 7'h20 == _myNewVec_80_T_3[6:0] ? myVec_32 : _GEN_6217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6219 = 7'h21 == _myNewVec_80_T_3[6:0] ? myVec_33 : _GEN_6218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6220 = 7'h22 == _myNewVec_80_T_3[6:0] ? myVec_34 : _GEN_6219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6221 = 7'h23 == _myNewVec_80_T_3[6:0] ? myVec_35 : _GEN_6220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6222 = 7'h24 == _myNewVec_80_T_3[6:0] ? myVec_36 : _GEN_6221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6223 = 7'h25 == _myNewVec_80_T_3[6:0] ? myVec_37 : _GEN_6222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6224 = 7'h26 == _myNewVec_80_T_3[6:0] ? myVec_38 : _GEN_6223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6225 = 7'h27 == _myNewVec_80_T_3[6:0] ? myVec_39 : _GEN_6224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6226 = 7'h28 == _myNewVec_80_T_3[6:0] ? myVec_40 : _GEN_6225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6227 = 7'h29 == _myNewVec_80_T_3[6:0] ? myVec_41 : _GEN_6226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6228 = 7'h2a == _myNewVec_80_T_3[6:0] ? myVec_42 : _GEN_6227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6229 = 7'h2b == _myNewVec_80_T_3[6:0] ? myVec_43 : _GEN_6228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6230 = 7'h2c == _myNewVec_80_T_3[6:0] ? myVec_44 : _GEN_6229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6231 = 7'h2d == _myNewVec_80_T_3[6:0] ? myVec_45 : _GEN_6230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6232 = 7'h2e == _myNewVec_80_T_3[6:0] ? myVec_46 : _GEN_6231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6233 = 7'h2f == _myNewVec_80_T_3[6:0] ? myVec_47 : _GEN_6232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6234 = 7'h30 == _myNewVec_80_T_3[6:0] ? myVec_48 : _GEN_6233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6235 = 7'h31 == _myNewVec_80_T_3[6:0] ? myVec_49 : _GEN_6234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6236 = 7'h32 == _myNewVec_80_T_3[6:0] ? myVec_50 : _GEN_6235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6237 = 7'h33 == _myNewVec_80_T_3[6:0] ? myVec_51 : _GEN_6236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6238 = 7'h34 == _myNewVec_80_T_3[6:0] ? myVec_52 : _GEN_6237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6239 = 7'h35 == _myNewVec_80_T_3[6:0] ? myVec_53 : _GEN_6238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6240 = 7'h36 == _myNewVec_80_T_3[6:0] ? myVec_54 : _GEN_6239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6241 = 7'h37 == _myNewVec_80_T_3[6:0] ? myVec_55 : _GEN_6240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6242 = 7'h38 == _myNewVec_80_T_3[6:0] ? myVec_56 : _GEN_6241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6243 = 7'h39 == _myNewVec_80_T_3[6:0] ? myVec_57 : _GEN_6242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6244 = 7'h3a == _myNewVec_80_T_3[6:0] ? myVec_58 : _GEN_6243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6245 = 7'h3b == _myNewVec_80_T_3[6:0] ? myVec_59 : _GEN_6244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6246 = 7'h3c == _myNewVec_80_T_3[6:0] ? myVec_60 : _GEN_6245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6247 = 7'h3d == _myNewVec_80_T_3[6:0] ? myVec_61 : _GEN_6246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6248 = 7'h3e == _myNewVec_80_T_3[6:0] ? myVec_62 : _GEN_6247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6249 = 7'h3f == _myNewVec_80_T_3[6:0] ? myVec_63 : _GEN_6248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6250 = 7'h40 == _myNewVec_80_T_3[6:0] ? myVec_64 : _GEN_6249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6251 = 7'h41 == _myNewVec_80_T_3[6:0] ? myVec_65 : _GEN_6250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6252 = 7'h42 == _myNewVec_80_T_3[6:0] ? myVec_66 : _GEN_6251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6253 = 7'h43 == _myNewVec_80_T_3[6:0] ? myVec_67 : _GEN_6252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6254 = 7'h44 == _myNewVec_80_T_3[6:0] ? myVec_68 : _GEN_6253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6255 = 7'h45 == _myNewVec_80_T_3[6:0] ? myVec_69 : _GEN_6254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6256 = 7'h46 == _myNewVec_80_T_3[6:0] ? myVec_70 : _GEN_6255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6257 = 7'h47 == _myNewVec_80_T_3[6:0] ? myVec_71 : _GEN_6256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6258 = 7'h48 == _myNewVec_80_T_3[6:0] ? myVec_72 : _GEN_6257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6259 = 7'h49 == _myNewVec_80_T_3[6:0] ? myVec_73 : _GEN_6258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6260 = 7'h4a == _myNewVec_80_T_3[6:0] ? myVec_74 : _GEN_6259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6261 = 7'h4b == _myNewVec_80_T_3[6:0] ? myVec_75 : _GEN_6260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6262 = 7'h4c == _myNewVec_80_T_3[6:0] ? myVec_76 : _GEN_6261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6263 = 7'h4d == _myNewVec_80_T_3[6:0] ? myVec_77 : _GEN_6262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6264 = 7'h4e == _myNewVec_80_T_3[6:0] ? myVec_78 : _GEN_6263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6265 = 7'h4f == _myNewVec_80_T_3[6:0] ? myVec_79 : _GEN_6264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6266 = 7'h50 == _myNewVec_80_T_3[6:0] ? myVec_80 : _GEN_6265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6267 = 7'h51 == _myNewVec_80_T_3[6:0] ? myVec_81 : _GEN_6266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6268 = 7'h52 == _myNewVec_80_T_3[6:0] ? myVec_82 : _GEN_6267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6269 = 7'h53 == _myNewVec_80_T_3[6:0] ? myVec_83 : _GEN_6268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6270 = 7'h54 == _myNewVec_80_T_3[6:0] ? myVec_84 : _GEN_6269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6271 = 7'h55 == _myNewVec_80_T_3[6:0] ? myVec_85 : _GEN_6270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6272 = 7'h56 == _myNewVec_80_T_3[6:0] ? myVec_86 : _GEN_6271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6273 = 7'h57 == _myNewVec_80_T_3[6:0] ? myVec_87 : _GEN_6272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6274 = 7'h58 == _myNewVec_80_T_3[6:0] ? myVec_88 : _GEN_6273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6275 = 7'h59 == _myNewVec_80_T_3[6:0] ? myVec_89 : _GEN_6274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6276 = 7'h5a == _myNewVec_80_T_3[6:0] ? myVec_90 : _GEN_6275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6277 = 7'h5b == _myNewVec_80_T_3[6:0] ? myVec_91 : _GEN_6276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6278 = 7'h5c == _myNewVec_80_T_3[6:0] ? myVec_92 : _GEN_6277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6279 = 7'h5d == _myNewVec_80_T_3[6:0] ? myVec_93 : _GEN_6278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6280 = 7'h5e == _myNewVec_80_T_3[6:0] ? myVec_94 : _GEN_6279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6281 = 7'h5f == _myNewVec_80_T_3[6:0] ? myVec_95 : _GEN_6280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6282 = 7'h60 == _myNewVec_80_T_3[6:0] ? myVec_96 : _GEN_6281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6283 = 7'h61 == _myNewVec_80_T_3[6:0] ? myVec_97 : _GEN_6282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6284 = 7'h62 == _myNewVec_80_T_3[6:0] ? myVec_98 : _GEN_6283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6285 = 7'h63 == _myNewVec_80_T_3[6:0] ? myVec_99 : _GEN_6284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6286 = 7'h64 == _myNewVec_80_T_3[6:0] ? myVec_100 : _GEN_6285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6287 = 7'h65 == _myNewVec_80_T_3[6:0] ? myVec_101 : _GEN_6286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6288 = 7'h66 == _myNewVec_80_T_3[6:0] ? myVec_102 : _GEN_6287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6289 = 7'h67 == _myNewVec_80_T_3[6:0] ? myVec_103 : _GEN_6288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6290 = 7'h68 == _myNewVec_80_T_3[6:0] ? myVec_104 : _GEN_6289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6291 = 7'h69 == _myNewVec_80_T_3[6:0] ? myVec_105 : _GEN_6290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6292 = 7'h6a == _myNewVec_80_T_3[6:0] ? myVec_106 : _GEN_6291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6293 = 7'h6b == _myNewVec_80_T_3[6:0] ? myVec_107 : _GEN_6292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6294 = 7'h6c == _myNewVec_80_T_3[6:0] ? myVec_108 : _GEN_6293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6295 = 7'h6d == _myNewVec_80_T_3[6:0] ? myVec_109 : _GEN_6294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6296 = 7'h6e == _myNewVec_80_T_3[6:0] ? myVec_110 : _GEN_6295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6297 = 7'h6f == _myNewVec_80_T_3[6:0] ? myVec_111 : _GEN_6296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6298 = 7'h70 == _myNewVec_80_T_3[6:0] ? myVec_112 : _GEN_6297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6299 = 7'h71 == _myNewVec_80_T_3[6:0] ? myVec_113 : _GEN_6298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6300 = 7'h72 == _myNewVec_80_T_3[6:0] ? myVec_114 : _GEN_6299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6301 = 7'h73 == _myNewVec_80_T_3[6:0] ? myVec_115 : _GEN_6300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6302 = 7'h74 == _myNewVec_80_T_3[6:0] ? myVec_116 : _GEN_6301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6303 = 7'h75 == _myNewVec_80_T_3[6:0] ? myVec_117 : _GEN_6302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6304 = 7'h76 == _myNewVec_80_T_3[6:0] ? myVec_118 : _GEN_6303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6305 = 7'h77 == _myNewVec_80_T_3[6:0] ? myVec_119 : _GEN_6304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6306 = 7'h78 == _myNewVec_80_T_3[6:0] ? myVec_120 : _GEN_6305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6307 = 7'h79 == _myNewVec_80_T_3[6:0] ? myVec_121 : _GEN_6306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6308 = 7'h7a == _myNewVec_80_T_3[6:0] ? myVec_122 : _GEN_6307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6309 = 7'h7b == _myNewVec_80_T_3[6:0] ? myVec_123 : _GEN_6308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6310 = 7'h7c == _myNewVec_80_T_3[6:0] ? myVec_124 : _GEN_6309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6311 = 7'h7d == _myNewVec_80_T_3[6:0] ? myVec_125 : _GEN_6310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6312 = 7'h7e == _myNewVec_80_T_3[6:0] ? myVec_126 : _GEN_6311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_80 = 7'h7f == _myNewVec_80_T_3[6:0] ? myVec_127 : _GEN_6312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [255:0] myNewWire_hi_lo_hi_lo = {myNewVec_87,myNewVec_86,myNewVec_85,myNewVec_84,myNewVec_83,myNewVec_82,
    myNewVec_81,myNewVec_80}; // @[hh_datapath_chisel.scala 238:27]
  wire [15:0] _myNewVec_79_T_3 = _myNewVec_127_T_1 + 16'h30; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_6315 = 7'h1 == _myNewVec_79_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6316 = 7'h2 == _myNewVec_79_T_3[6:0] ? myVec_2 : _GEN_6315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6317 = 7'h3 == _myNewVec_79_T_3[6:0] ? myVec_3 : _GEN_6316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6318 = 7'h4 == _myNewVec_79_T_3[6:0] ? myVec_4 : _GEN_6317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6319 = 7'h5 == _myNewVec_79_T_3[6:0] ? myVec_5 : _GEN_6318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6320 = 7'h6 == _myNewVec_79_T_3[6:0] ? myVec_6 : _GEN_6319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6321 = 7'h7 == _myNewVec_79_T_3[6:0] ? myVec_7 : _GEN_6320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6322 = 7'h8 == _myNewVec_79_T_3[6:0] ? myVec_8 : _GEN_6321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6323 = 7'h9 == _myNewVec_79_T_3[6:0] ? myVec_9 : _GEN_6322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6324 = 7'ha == _myNewVec_79_T_3[6:0] ? myVec_10 : _GEN_6323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6325 = 7'hb == _myNewVec_79_T_3[6:0] ? myVec_11 : _GEN_6324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6326 = 7'hc == _myNewVec_79_T_3[6:0] ? myVec_12 : _GEN_6325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6327 = 7'hd == _myNewVec_79_T_3[6:0] ? myVec_13 : _GEN_6326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6328 = 7'he == _myNewVec_79_T_3[6:0] ? myVec_14 : _GEN_6327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6329 = 7'hf == _myNewVec_79_T_3[6:0] ? myVec_15 : _GEN_6328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6330 = 7'h10 == _myNewVec_79_T_3[6:0] ? myVec_16 : _GEN_6329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6331 = 7'h11 == _myNewVec_79_T_3[6:0] ? myVec_17 : _GEN_6330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6332 = 7'h12 == _myNewVec_79_T_3[6:0] ? myVec_18 : _GEN_6331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6333 = 7'h13 == _myNewVec_79_T_3[6:0] ? myVec_19 : _GEN_6332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6334 = 7'h14 == _myNewVec_79_T_3[6:0] ? myVec_20 : _GEN_6333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6335 = 7'h15 == _myNewVec_79_T_3[6:0] ? myVec_21 : _GEN_6334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6336 = 7'h16 == _myNewVec_79_T_3[6:0] ? myVec_22 : _GEN_6335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6337 = 7'h17 == _myNewVec_79_T_3[6:0] ? myVec_23 : _GEN_6336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6338 = 7'h18 == _myNewVec_79_T_3[6:0] ? myVec_24 : _GEN_6337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6339 = 7'h19 == _myNewVec_79_T_3[6:0] ? myVec_25 : _GEN_6338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6340 = 7'h1a == _myNewVec_79_T_3[6:0] ? myVec_26 : _GEN_6339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6341 = 7'h1b == _myNewVec_79_T_3[6:0] ? myVec_27 : _GEN_6340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6342 = 7'h1c == _myNewVec_79_T_3[6:0] ? myVec_28 : _GEN_6341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6343 = 7'h1d == _myNewVec_79_T_3[6:0] ? myVec_29 : _GEN_6342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6344 = 7'h1e == _myNewVec_79_T_3[6:0] ? myVec_30 : _GEN_6343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6345 = 7'h1f == _myNewVec_79_T_3[6:0] ? myVec_31 : _GEN_6344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6346 = 7'h20 == _myNewVec_79_T_3[6:0] ? myVec_32 : _GEN_6345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6347 = 7'h21 == _myNewVec_79_T_3[6:0] ? myVec_33 : _GEN_6346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6348 = 7'h22 == _myNewVec_79_T_3[6:0] ? myVec_34 : _GEN_6347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6349 = 7'h23 == _myNewVec_79_T_3[6:0] ? myVec_35 : _GEN_6348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6350 = 7'h24 == _myNewVec_79_T_3[6:0] ? myVec_36 : _GEN_6349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6351 = 7'h25 == _myNewVec_79_T_3[6:0] ? myVec_37 : _GEN_6350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6352 = 7'h26 == _myNewVec_79_T_3[6:0] ? myVec_38 : _GEN_6351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6353 = 7'h27 == _myNewVec_79_T_3[6:0] ? myVec_39 : _GEN_6352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6354 = 7'h28 == _myNewVec_79_T_3[6:0] ? myVec_40 : _GEN_6353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6355 = 7'h29 == _myNewVec_79_T_3[6:0] ? myVec_41 : _GEN_6354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6356 = 7'h2a == _myNewVec_79_T_3[6:0] ? myVec_42 : _GEN_6355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6357 = 7'h2b == _myNewVec_79_T_3[6:0] ? myVec_43 : _GEN_6356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6358 = 7'h2c == _myNewVec_79_T_3[6:0] ? myVec_44 : _GEN_6357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6359 = 7'h2d == _myNewVec_79_T_3[6:0] ? myVec_45 : _GEN_6358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6360 = 7'h2e == _myNewVec_79_T_3[6:0] ? myVec_46 : _GEN_6359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6361 = 7'h2f == _myNewVec_79_T_3[6:0] ? myVec_47 : _GEN_6360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6362 = 7'h30 == _myNewVec_79_T_3[6:0] ? myVec_48 : _GEN_6361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6363 = 7'h31 == _myNewVec_79_T_3[6:0] ? myVec_49 : _GEN_6362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6364 = 7'h32 == _myNewVec_79_T_3[6:0] ? myVec_50 : _GEN_6363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6365 = 7'h33 == _myNewVec_79_T_3[6:0] ? myVec_51 : _GEN_6364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6366 = 7'h34 == _myNewVec_79_T_3[6:0] ? myVec_52 : _GEN_6365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6367 = 7'h35 == _myNewVec_79_T_3[6:0] ? myVec_53 : _GEN_6366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6368 = 7'h36 == _myNewVec_79_T_3[6:0] ? myVec_54 : _GEN_6367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6369 = 7'h37 == _myNewVec_79_T_3[6:0] ? myVec_55 : _GEN_6368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6370 = 7'h38 == _myNewVec_79_T_3[6:0] ? myVec_56 : _GEN_6369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6371 = 7'h39 == _myNewVec_79_T_3[6:0] ? myVec_57 : _GEN_6370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6372 = 7'h3a == _myNewVec_79_T_3[6:0] ? myVec_58 : _GEN_6371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6373 = 7'h3b == _myNewVec_79_T_3[6:0] ? myVec_59 : _GEN_6372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6374 = 7'h3c == _myNewVec_79_T_3[6:0] ? myVec_60 : _GEN_6373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6375 = 7'h3d == _myNewVec_79_T_3[6:0] ? myVec_61 : _GEN_6374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6376 = 7'h3e == _myNewVec_79_T_3[6:0] ? myVec_62 : _GEN_6375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6377 = 7'h3f == _myNewVec_79_T_3[6:0] ? myVec_63 : _GEN_6376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6378 = 7'h40 == _myNewVec_79_T_3[6:0] ? myVec_64 : _GEN_6377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6379 = 7'h41 == _myNewVec_79_T_3[6:0] ? myVec_65 : _GEN_6378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6380 = 7'h42 == _myNewVec_79_T_3[6:0] ? myVec_66 : _GEN_6379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6381 = 7'h43 == _myNewVec_79_T_3[6:0] ? myVec_67 : _GEN_6380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6382 = 7'h44 == _myNewVec_79_T_3[6:0] ? myVec_68 : _GEN_6381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6383 = 7'h45 == _myNewVec_79_T_3[6:0] ? myVec_69 : _GEN_6382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6384 = 7'h46 == _myNewVec_79_T_3[6:0] ? myVec_70 : _GEN_6383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6385 = 7'h47 == _myNewVec_79_T_3[6:0] ? myVec_71 : _GEN_6384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6386 = 7'h48 == _myNewVec_79_T_3[6:0] ? myVec_72 : _GEN_6385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6387 = 7'h49 == _myNewVec_79_T_3[6:0] ? myVec_73 : _GEN_6386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6388 = 7'h4a == _myNewVec_79_T_3[6:0] ? myVec_74 : _GEN_6387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6389 = 7'h4b == _myNewVec_79_T_3[6:0] ? myVec_75 : _GEN_6388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6390 = 7'h4c == _myNewVec_79_T_3[6:0] ? myVec_76 : _GEN_6389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6391 = 7'h4d == _myNewVec_79_T_3[6:0] ? myVec_77 : _GEN_6390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6392 = 7'h4e == _myNewVec_79_T_3[6:0] ? myVec_78 : _GEN_6391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6393 = 7'h4f == _myNewVec_79_T_3[6:0] ? myVec_79 : _GEN_6392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6394 = 7'h50 == _myNewVec_79_T_3[6:0] ? myVec_80 : _GEN_6393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6395 = 7'h51 == _myNewVec_79_T_3[6:0] ? myVec_81 : _GEN_6394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6396 = 7'h52 == _myNewVec_79_T_3[6:0] ? myVec_82 : _GEN_6395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6397 = 7'h53 == _myNewVec_79_T_3[6:0] ? myVec_83 : _GEN_6396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6398 = 7'h54 == _myNewVec_79_T_3[6:0] ? myVec_84 : _GEN_6397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6399 = 7'h55 == _myNewVec_79_T_3[6:0] ? myVec_85 : _GEN_6398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6400 = 7'h56 == _myNewVec_79_T_3[6:0] ? myVec_86 : _GEN_6399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6401 = 7'h57 == _myNewVec_79_T_3[6:0] ? myVec_87 : _GEN_6400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6402 = 7'h58 == _myNewVec_79_T_3[6:0] ? myVec_88 : _GEN_6401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6403 = 7'h59 == _myNewVec_79_T_3[6:0] ? myVec_89 : _GEN_6402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6404 = 7'h5a == _myNewVec_79_T_3[6:0] ? myVec_90 : _GEN_6403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6405 = 7'h5b == _myNewVec_79_T_3[6:0] ? myVec_91 : _GEN_6404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6406 = 7'h5c == _myNewVec_79_T_3[6:0] ? myVec_92 : _GEN_6405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6407 = 7'h5d == _myNewVec_79_T_3[6:0] ? myVec_93 : _GEN_6406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6408 = 7'h5e == _myNewVec_79_T_3[6:0] ? myVec_94 : _GEN_6407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6409 = 7'h5f == _myNewVec_79_T_3[6:0] ? myVec_95 : _GEN_6408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6410 = 7'h60 == _myNewVec_79_T_3[6:0] ? myVec_96 : _GEN_6409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6411 = 7'h61 == _myNewVec_79_T_3[6:0] ? myVec_97 : _GEN_6410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6412 = 7'h62 == _myNewVec_79_T_3[6:0] ? myVec_98 : _GEN_6411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6413 = 7'h63 == _myNewVec_79_T_3[6:0] ? myVec_99 : _GEN_6412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6414 = 7'h64 == _myNewVec_79_T_3[6:0] ? myVec_100 : _GEN_6413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6415 = 7'h65 == _myNewVec_79_T_3[6:0] ? myVec_101 : _GEN_6414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6416 = 7'h66 == _myNewVec_79_T_3[6:0] ? myVec_102 : _GEN_6415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6417 = 7'h67 == _myNewVec_79_T_3[6:0] ? myVec_103 : _GEN_6416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6418 = 7'h68 == _myNewVec_79_T_3[6:0] ? myVec_104 : _GEN_6417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6419 = 7'h69 == _myNewVec_79_T_3[6:0] ? myVec_105 : _GEN_6418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6420 = 7'h6a == _myNewVec_79_T_3[6:0] ? myVec_106 : _GEN_6419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6421 = 7'h6b == _myNewVec_79_T_3[6:0] ? myVec_107 : _GEN_6420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6422 = 7'h6c == _myNewVec_79_T_3[6:0] ? myVec_108 : _GEN_6421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6423 = 7'h6d == _myNewVec_79_T_3[6:0] ? myVec_109 : _GEN_6422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6424 = 7'h6e == _myNewVec_79_T_3[6:0] ? myVec_110 : _GEN_6423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6425 = 7'h6f == _myNewVec_79_T_3[6:0] ? myVec_111 : _GEN_6424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6426 = 7'h70 == _myNewVec_79_T_3[6:0] ? myVec_112 : _GEN_6425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6427 = 7'h71 == _myNewVec_79_T_3[6:0] ? myVec_113 : _GEN_6426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6428 = 7'h72 == _myNewVec_79_T_3[6:0] ? myVec_114 : _GEN_6427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6429 = 7'h73 == _myNewVec_79_T_3[6:0] ? myVec_115 : _GEN_6428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6430 = 7'h74 == _myNewVec_79_T_3[6:0] ? myVec_116 : _GEN_6429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6431 = 7'h75 == _myNewVec_79_T_3[6:0] ? myVec_117 : _GEN_6430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6432 = 7'h76 == _myNewVec_79_T_3[6:0] ? myVec_118 : _GEN_6431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6433 = 7'h77 == _myNewVec_79_T_3[6:0] ? myVec_119 : _GEN_6432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6434 = 7'h78 == _myNewVec_79_T_3[6:0] ? myVec_120 : _GEN_6433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6435 = 7'h79 == _myNewVec_79_T_3[6:0] ? myVec_121 : _GEN_6434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6436 = 7'h7a == _myNewVec_79_T_3[6:0] ? myVec_122 : _GEN_6435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6437 = 7'h7b == _myNewVec_79_T_3[6:0] ? myVec_123 : _GEN_6436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6438 = 7'h7c == _myNewVec_79_T_3[6:0] ? myVec_124 : _GEN_6437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6439 = 7'h7d == _myNewVec_79_T_3[6:0] ? myVec_125 : _GEN_6438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6440 = 7'h7e == _myNewVec_79_T_3[6:0] ? myVec_126 : _GEN_6439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_79 = 7'h7f == _myNewVec_79_T_3[6:0] ? myVec_127 : _GEN_6440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_78_T_3 = _myNewVec_127_T_1 + 16'h31; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_6443 = 7'h1 == _myNewVec_78_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6444 = 7'h2 == _myNewVec_78_T_3[6:0] ? myVec_2 : _GEN_6443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6445 = 7'h3 == _myNewVec_78_T_3[6:0] ? myVec_3 : _GEN_6444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6446 = 7'h4 == _myNewVec_78_T_3[6:0] ? myVec_4 : _GEN_6445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6447 = 7'h5 == _myNewVec_78_T_3[6:0] ? myVec_5 : _GEN_6446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6448 = 7'h6 == _myNewVec_78_T_3[6:0] ? myVec_6 : _GEN_6447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6449 = 7'h7 == _myNewVec_78_T_3[6:0] ? myVec_7 : _GEN_6448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6450 = 7'h8 == _myNewVec_78_T_3[6:0] ? myVec_8 : _GEN_6449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6451 = 7'h9 == _myNewVec_78_T_3[6:0] ? myVec_9 : _GEN_6450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6452 = 7'ha == _myNewVec_78_T_3[6:0] ? myVec_10 : _GEN_6451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6453 = 7'hb == _myNewVec_78_T_3[6:0] ? myVec_11 : _GEN_6452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6454 = 7'hc == _myNewVec_78_T_3[6:0] ? myVec_12 : _GEN_6453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6455 = 7'hd == _myNewVec_78_T_3[6:0] ? myVec_13 : _GEN_6454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6456 = 7'he == _myNewVec_78_T_3[6:0] ? myVec_14 : _GEN_6455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6457 = 7'hf == _myNewVec_78_T_3[6:0] ? myVec_15 : _GEN_6456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6458 = 7'h10 == _myNewVec_78_T_3[6:0] ? myVec_16 : _GEN_6457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6459 = 7'h11 == _myNewVec_78_T_3[6:0] ? myVec_17 : _GEN_6458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6460 = 7'h12 == _myNewVec_78_T_3[6:0] ? myVec_18 : _GEN_6459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6461 = 7'h13 == _myNewVec_78_T_3[6:0] ? myVec_19 : _GEN_6460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6462 = 7'h14 == _myNewVec_78_T_3[6:0] ? myVec_20 : _GEN_6461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6463 = 7'h15 == _myNewVec_78_T_3[6:0] ? myVec_21 : _GEN_6462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6464 = 7'h16 == _myNewVec_78_T_3[6:0] ? myVec_22 : _GEN_6463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6465 = 7'h17 == _myNewVec_78_T_3[6:0] ? myVec_23 : _GEN_6464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6466 = 7'h18 == _myNewVec_78_T_3[6:0] ? myVec_24 : _GEN_6465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6467 = 7'h19 == _myNewVec_78_T_3[6:0] ? myVec_25 : _GEN_6466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6468 = 7'h1a == _myNewVec_78_T_3[6:0] ? myVec_26 : _GEN_6467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6469 = 7'h1b == _myNewVec_78_T_3[6:0] ? myVec_27 : _GEN_6468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6470 = 7'h1c == _myNewVec_78_T_3[6:0] ? myVec_28 : _GEN_6469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6471 = 7'h1d == _myNewVec_78_T_3[6:0] ? myVec_29 : _GEN_6470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6472 = 7'h1e == _myNewVec_78_T_3[6:0] ? myVec_30 : _GEN_6471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6473 = 7'h1f == _myNewVec_78_T_3[6:0] ? myVec_31 : _GEN_6472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6474 = 7'h20 == _myNewVec_78_T_3[6:0] ? myVec_32 : _GEN_6473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6475 = 7'h21 == _myNewVec_78_T_3[6:0] ? myVec_33 : _GEN_6474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6476 = 7'h22 == _myNewVec_78_T_3[6:0] ? myVec_34 : _GEN_6475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6477 = 7'h23 == _myNewVec_78_T_3[6:0] ? myVec_35 : _GEN_6476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6478 = 7'h24 == _myNewVec_78_T_3[6:0] ? myVec_36 : _GEN_6477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6479 = 7'h25 == _myNewVec_78_T_3[6:0] ? myVec_37 : _GEN_6478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6480 = 7'h26 == _myNewVec_78_T_3[6:0] ? myVec_38 : _GEN_6479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6481 = 7'h27 == _myNewVec_78_T_3[6:0] ? myVec_39 : _GEN_6480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6482 = 7'h28 == _myNewVec_78_T_3[6:0] ? myVec_40 : _GEN_6481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6483 = 7'h29 == _myNewVec_78_T_3[6:0] ? myVec_41 : _GEN_6482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6484 = 7'h2a == _myNewVec_78_T_3[6:0] ? myVec_42 : _GEN_6483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6485 = 7'h2b == _myNewVec_78_T_3[6:0] ? myVec_43 : _GEN_6484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6486 = 7'h2c == _myNewVec_78_T_3[6:0] ? myVec_44 : _GEN_6485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6487 = 7'h2d == _myNewVec_78_T_3[6:0] ? myVec_45 : _GEN_6486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6488 = 7'h2e == _myNewVec_78_T_3[6:0] ? myVec_46 : _GEN_6487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6489 = 7'h2f == _myNewVec_78_T_3[6:0] ? myVec_47 : _GEN_6488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6490 = 7'h30 == _myNewVec_78_T_3[6:0] ? myVec_48 : _GEN_6489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6491 = 7'h31 == _myNewVec_78_T_3[6:0] ? myVec_49 : _GEN_6490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6492 = 7'h32 == _myNewVec_78_T_3[6:0] ? myVec_50 : _GEN_6491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6493 = 7'h33 == _myNewVec_78_T_3[6:0] ? myVec_51 : _GEN_6492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6494 = 7'h34 == _myNewVec_78_T_3[6:0] ? myVec_52 : _GEN_6493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6495 = 7'h35 == _myNewVec_78_T_3[6:0] ? myVec_53 : _GEN_6494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6496 = 7'h36 == _myNewVec_78_T_3[6:0] ? myVec_54 : _GEN_6495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6497 = 7'h37 == _myNewVec_78_T_3[6:0] ? myVec_55 : _GEN_6496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6498 = 7'h38 == _myNewVec_78_T_3[6:0] ? myVec_56 : _GEN_6497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6499 = 7'h39 == _myNewVec_78_T_3[6:0] ? myVec_57 : _GEN_6498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6500 = 7'h3a == _myNewVec_78_T_3[6:0] ? myVec_58 : _GEN_6499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6501 = 7'h3b == _myNewVec_78_T_3[6:0] ? myVec_59 : _GEN_6500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6502 = 7'h3c == _myNewVec_78_T_3[6:0] ? myVec_60 : _GEN_6501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6503 = 7'h3d == _myNewVec_78_T_3[6:0] ? myVec_61 : _GEN_6502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6504 = 7'h3e == _myNewVec_78_T_3[6:0] ? myVec_62 : _GEN_6503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6505 = 7'h3f == _myNewVec_78_T_3[6:0] ? myVec_63 : _GEN_6504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6506 = 7'h40 == _myNewVec_78_T_3[6:0] ? myVec_64 : _GEN_6505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6507 = 7'h41 == _myNewVec_78_T_3[6:0] ? myVec_65 : _GEN_6506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6508 = 7'h42 == _myNewVec_78_T_3[6:0] ? myVec_66 : _GEN_6507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6509 = 7'h43 == _myNewVec_78_T_3[6:0] ? myVec_67 : _GEN_6508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6510 = 7'h44 == _myNewVec_78_T_3[6:0] ? myVec_68 : _GEN_6509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6511 = 7'h45 == _myNewVec_78_T_3[6:0] ? myVec_69 : _GEN_6510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6512 = 7'h46 == _myNewVec_78_T_3[6:0] ? myVec_70 : _GEN_6511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6513 = 7'h47 == _myNewVec_78_T_3[6:0] ? myVec_71 : _GEN_6512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6514 = 7'h48 == _myNewVec_78_T_3[6:0] ? myVec_72 : _GEN_6513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6515 = 7'h49 == _myNewVec_78_T_3[6:0] ? myVec_73 : _GEN_6514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6516 = 7'h4a == _myNewVec_78_T_3[6:0] ? myVec_74 : _GEN_6515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6517 = 7'h4b == _myNewVec_78_T_3[6:0] ? myVec_75 : _GEN_6516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6518 = 7'h4c == _myNewVec_78_T_3[6:0] ? myVec_76 : _GEN_6517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6519 = 7'h4d == _myNewVec_78_T_3[6:0] ? myVec_77 : _GEN_6518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6520 = 7'h4e == _myNewVec_78_T_3[6:0] ? myVec_78 : _GEN_6519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6521 = 7'h4f == _myNewVec_78_T_3[6:0] ? myVec_79 : _GEN_6520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6522 = 7'h50 == _myNewVec_78_T_3[6:0] ? myVec_80 : _GEN_6521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6523 = 7'h51 == _myNewVec_78_T_3[6:0] ? myVec_81 : _GEN_6522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6524 = 7'h52 == _myNewVec_78_T_3[6:0] ? myVec_82 : _GEN_6523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6525 = 7'h53 == _myNewVec_78_T_3[6:0] ? myVec_83 : _GEN_6524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6526 = 7'h54 == _myNewVec_78_T_3[6:0] ? myVec_84 : _GEN_6525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6527 = 7'h55 == _myNewVec_78_T_3[6:0] ? myVec_85 : _GEN_6526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6528 = 7'h56 == _myNewVec_78_T_3[6:0] ? myVec_86 : _GEN_6527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6529 = 7'h57 == _myNewVec_78_T_3[6:0] ? myVec_87 : _GEN_6528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6530 = 7'h58 == _myNewVec_78_T_3[6:0] ? myVec_88 : _GEN_6529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6531 = 7'h59 == _myNewVec_78_T_3[6:0] ? myVec_89 : _GEN_6530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6532 = 7'h5a == _myNewVec_78_T_3[6:0] ? myVec_90 : _GEN_6531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6533 = 7'h5b == _myNewVec_78_T_3[6:0] ? myVec_91 : _GEN_6532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6534 = 7'h5c == _myNewVec_78_T_3[6:0] ? myVec_92 : _GEN_6533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6535 = 7'h5d == _myNewVec_78_T_3[6:0] ? myVec_93 : _GEN_6534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6536 = 7'h5e == _myNewVec_78_T_3[6:0] ? myVec_94 : _GEN_6535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6537 = 7'h5f == _myNewVec_78_T_3[6:0] ? myVec_95 : _GEN_6536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6538 = 7'h60 == _myNewVec_78_T_3[6:0] ? myVec_96 : _GEN_6537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6539 = 7'h61 == _myNewVec_78_T_3[6:0] ? myVec_97 : _GEN_6538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6540 = 7'h62 == _myNewVec_78_T_3[6:0] ? myVec_98 : _GEN_6539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6541 = 7'h63 == _myNewVec_78_T_3[6:0] ? myVec_99 : _GEN_6540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6542 = 7'h64 == _myNewVec_78_T_3[6:0] ? myVec_100 : _GEN_6541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6543 = 7'h65 == _myNewVec_78_T_3[6:0] ? myVec_101 : _GEN_6542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6544 = 7'h66 == _myNewVec_78_T_3[6:0] ? myVec_102 : _GEN_6543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6545 = 7'h67 == _myNewVec_78_T_3[6:0] ? myVec_103 : _GEN_6544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6546 = 7'h68 == _myNewVec_78_T_3[6:0] ? myVec_104 : _GEN_6545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6547 = 7'h69 == _myNewVec_78_T_3[6:0] ? myVec_105 : _GEN_6546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6548 = 7'h6a == _myNewVec_78_T_3[6:0] ? myVec_106 : _GEN_6547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6549 = 7'h6b == _myNewVec_78_T_3[6:0] ? myVec_107 : _GEN_6548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6550 = 7'h6c == _myNewVec_78_T_3[6:0] ? myVec_108 : _GEN_6549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6551 = 7'h6d == _myNewVec_78_T_3[6:0] ? myVec_109 : _GEN_6550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6552 = 7'h6e == _myNewVec_78_T_3[6:0] ? myVec_110 : _GEN_6551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6553 = 7'h6f == _myNewVec_78_T_3[6:0] ? myVec_111 : _GEN_6552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6554 = 7'h70 == _myNewVec_78_T_3[6:0] ? myVec_112 : _GEN_6553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6555 = 7'h71 == _myNewVec_78_T_3[6:0] ? myVec_113 : _GEN_6554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6556 = 7'h72 == _myNewVec_78_T_3[6:0] ? myVec_114 : _GEN_6555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6557 = 7'h73 == _myNewVec_78_T_3[6:0] ? myVec_115 : _GEN_6556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6558 = 7'h74 == _myNewVec_78_T_3[6:0] ? myVec_116 : _GEN_6557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6559 = 7'h75 == _myNewVec_78_T_3[6:0] ? myVec_117 : _GEN_6558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6560 = 7'h76 == _myNewVec_78_T_3[6:0] ? myVec_118 : _GEN_6559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6561 = 7'h77 == _myNewVec_78_T_3[6:0] ? myVec_119 : _GEN_6560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6562 = 7'h78 == _myNewVec_78_T_3[6:0] ? myVec_120 : _GEN_6561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6563 = 7'h79 == _myNewVec_78_T_3[6:0] ? myVec_121 : _GEN_6562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6564 = 7'h7a == _myNewVec_78_T_3[6:0] ? myVec_122 : _GEN_6563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6565 = 7'h7b == _myNewVec_78_T_3[6:0] ? myVec_123 : _GEN_6564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6566 = 7'h7c == _myNewVec_78_T_3[6:0] ? myVec_124 : _GEN_6565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6567 = 7'h7d == _myNewVec_78_T_3[6:0] ? myVec_125 : _GEN_6566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6568 = 7'h7e == _myNewVec_78_T_3[6:0] ? myVec_126 : _GEN_6567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_78 = 7'h7f == _myNewVec_78_T_3[6:0] ? myVec_127 : _GEN_6568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_77_T_3 = _myNewVec_127_T_1 + 16'h32; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_6571 = 7'h1 == _myNewVec_77_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6572 = 7'h2 == _myNewVec_77_T_3[6:0] ? myVec_2 : _GEN_6571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6573 = 7'h3 == _myNewVec_77_T_3[6:0] ? myVec_3 : _GEN_6572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6574 = 7'h4 == _myNewVec_77_T_3[6:0] ? myVec_4 : _GEN_6573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6575 = 7'h5 == _myNewVec_77_T_3[6:0] ? myVec_5 : _GEN_6574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6576 = 7'h6 == _myNewVec_77_T_3[6:0] ? myVec_6 : _GEN_6575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6577 = 7'h7 == _myNewVec_77_T_3[6:0] ? myVec_7 : _GEN_6576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6578 = 7'h8 == _myNewVec_77_T_3[6:0] ? myVec_8 : _GEN_6577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6579 = 7'h9 == _myNewVec_77_T_3[6:0] ? myVec_9 : _GEN_6578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6580 = 7'ha == _myNewVec_77_T_3[6:0] ? myVec_10 : _GEN_6579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6581 = 7'hb == _myNewVec_77_T_3[6:0] ? myVec_11 : _GEN_6580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6582 = 7'hc == _myNewVec_77_T_3[6:0] ? myVec_12 : _GEN_6581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6583 = 7'hd == _myNewVec_77_T_3[6:0] ? myVec_13 : _GEN_6582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6584 = 7'he == _myNewVec_77_T_3[6:0] ? myVec_14 : _GEN_6583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6585 = 7'hf == _myNewVec_77_T_3[6:0] ? myVec_15 : _GEN_6584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6586 = 7'h10 == _myNewVec_77_T_3[6:0] ? myVec_16 : _GEN_6585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6587 = 7'h11 == _myNewVec_77_T_3[6:0] ? myVec_17 : _GEN_6586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6588 = 7'h12 == _myNewVec_77_T_3[6:0] ? myVec_18 : _GEN_6587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6589 = 7'h13 == _myNewVec_77_T_3[6:0] ? myVec_19 : _GEN_6588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6590 = 7'h14 == _myNewVec_77_T_3[6:0] ? myVec_20 : _GEN_6589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6591 = 7'h15 == _myNewVec_77_T_3[6:0] ? myVec_21 : _GEN_6590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6592 = 7'h16 == _myNewVec_77_T_3[6:0] ? myVec_22 : _GEN_6591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6593 = 7'h17 == _myNewVec_77_T_3[6:0] ? myVec_23 : _GEN_6592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6594 = 7'h18 == _myNewVec_77_T_3[6:0] ? myVec_24 : _GEN_6593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6595 = 7'h19 == _myNewVec_77_T_3[6:0] ? myVec_25 : _GEN_6594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6596 = 7'h1a == _myNewVec_77_T_3[6:0] ? myVec_26 : _GEN_6595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6597 = 7'h1b == _myNewVec_77_T_3[6:0] ? myVec_27 : _GEN_6596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6598 = 7'h1c == _myNewVec_77_T_3[6:0] ? myVec_28 : _GEN_6597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6599 = 7'h1d == _myNewVec_77_T_3[6:0] ? myVec_29 : _GEN_6598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6600 = 7'h1e == _myNewVec_77_T_3[6:0] ? myVec_30 : _GEN_6599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6601 = 7'h1f == _myNewVec_77_T_3[6:0] ? myVec_31 : _GEN_6600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6602 = 7'h20 == _myNewVec_77_T_3[6:0] ? myVec_32 : _GEN_6601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6603 = 7'h21 == _myNewVec_77_T_3[6:0] ? myVec_33 : _GEN_6602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6604 = 7'h22 == _myNewVec_77_T_3[6:0] ? myVec_34 : _GEN_6603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6605 = 7'h23 == _myNewVec_77_T_3[6:0] ? myVec_35 : _GEN_6604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6606 = 7'h24 == _myNewVec_77_T_3[6:0] ? myVec_36 : _GEN_6605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6607 = 7'h25 == _myNewVec_77_T_3[6:0] ? myVec_37 : _GEN_6606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6608 = 7'h26 == _myNewVec_77_T_3[6:0] ? myVec_38 : _GEN_6607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6609 = 7'h27 == _myNewVec_77_T_3[6:0] ? myVec_39 : _GEN_6608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6610 = 7'h28 == _myNewVec_77_T_3[6:0] ? myVec_40 : _GEN_6609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6611 = 7'h29 == _myNewVec_77_T_3[6:0] ? myVec_41 : _GEN_6610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6612 = 7'h2a == _myNewVec_77_T_3[6:0] ? myVec_42 : _GEN_6611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6613 = 7'h2b == _myNewVec_77_T_3[6:0] ? myVec_43 : _GEN_6612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6614 = 7'h2c == _myNewVec_77_T_3[6:0] ? myVec_44 : _GEN_6613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6615 = 7'h2d == _myNewVec_77_T_3[6:0] ? myVec_45 : _GEN_6614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6616 = 7'h2e == _myNewVec_77_T_3[6:0] ? myVec_46 : _GEN_6615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6617 = 7'h2f == _myNewVec_77_T_3[6:0] ? myVec_47 : _GEN_6616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6618 = 7'h30 == _myNewVec_77_T_3[6:0] ? myVec_48 : _GEN_6617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6619 = 7'h31 == _myNewVec_77_T_3[6:0] ? myVec_49 : _GEN_6618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6620 = 7'h32 == _myNewVec_77_T_3[6:0] ? myVec_50 : _GEN_6619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6621 = 7'h33 == _myNewVec_77_T_3[6:0] ? myVec_51 : _GEN_6620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6622 = 7'h34 == _myNewVec_77_T_3[6:0] ? myVec_52 : _GEN_6621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6623 = 7'h35 == _myNewVec_77_T_3[6:0] ? myVec_53 : _GEN_6622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6624 = 7'h36 == _myNewVec_77_T_3[6:0] ? myVec_54 : _GEN_6623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6625 = 7'h37 == _myNewVec_77_T_3[6:0] ? myVec_55 : _GEN_6624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6626 = 7'h38 == _myNewVec_77_T_3[6:0] ? myVec_56 : _GEN_6625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6627 = 7'h39 == _myNewVec_77_T_3[6:0] ? myVec_57 : _GEN_6626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6628 = 7'h3a == _myNewVec_77_T_3[6:0] ? myVec_58 : _GEN_6627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6629 = 7'h3b == _myNewVec_77_T_3[6:0] ? myVec_59 : _GEN_6628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6630 = 7'h3c == _myNewVec_77_T_3[6:0] ? myVec_60 : _GEN_6629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6631 = 7'h3d == _myNewVec_77_T_3[6:0] ? myVec_61 : _GEN_6630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6632 = 7'h3e == _myNewVec_77_T_3[6:0] ? myVec_62 : _GEN_6631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6633 = 7'h3f == _myNewVec_77_T_3[6:0] ? myVec_63 : _GEN_6632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6634 = 7'h40 == _myNewVec_77_T_3[6:0] ? myVec_64 : _GEN_6633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6635 = 7'h41 == _myNewVec_77_T_3[6:0] ? myVec_65 : _GEN_6634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6636 = 7'h42 == _myNewVec_77_T_3[6:0] ? myVec_66 : _GEN_6635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6637 = 7'h43 == _myNewVec_77_T_3[6:0] ? myVec_67 : _GEN_6636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6638 = 7'h44 == _myNewVec_77_T_3[6:0] ? myVec_68 : _GEN_6637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6639 = 7'h45 == _myNewVec_77_T_3[6:0] ? myVec_69 : _GEN_6638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6640 = 7'h46 == _myNewVec_77_T_3[6:0] ? myVec_70 : _GEN_6639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6641 = 7'h47 == _myNewVec_77_T_3[6:0] ? myVec_71 : _GEN_6640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6642 = 7'h48 == _myNewVec_77_T_3[6:0] ? myVec_72 : _GEN_6641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6643 = 7'h49 == _myNewVec_77_T_3[6:0] ? myVec_73 : _GEN_6642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6644 = 7'h4a == _myNewVec_77_T_3[6:0] ? myVec_74 : _GEN_6643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6645 = 7'h4b == _myNewVec_77_T_3[6:0] ? myVec_75 : _GEN_6644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6646 = 7'h4c == _myNewVec_77_T_3[6:0] ? myVec_76 : _GEN_6645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6647 = 7'h4d == _myNewVec_77_T_3[6:0] ? myVec_77 : _GEN_6646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6648 = 7'h4e == _myNewVec_77_T_3[6:0] ? myVec_78 : _GEN_6647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6649 = 7'h4f == _myNewVec_77_T_3[6:0] ? myVec_79 : _GEN_6648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6650 = 7'h50 == _myNewVec_77_T_3[6:0] ? myVec_80 : _GEN_6649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6651 = 7'h51 == _myNewVec_77_T_3[6:0] ? myVec_81 : _GEN_6650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6652 = 7'h52 == _myNewVec_77_T_3[6:0] ? myVec_82 : _GEN_6651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6653 = 7'h53 == _myNewVec_77_T_3[6:0] ? myVec_83 : _GEN_6652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6654 = 7'h54 == _myNewVec_77_T_3[6:0] ? myVec_84 : _GEN_6653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6655 = 7'h55 == _myNewVec_77_T_3[6:0] ? myVec_85 : _GEN_6654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6656 = 7'h56 == _myNewVec_77_T_3[6:0] ? myVec_86 : _GEN_6655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6657 = 7'h57 == _myNewVec_77_T_3[6:0] ? myVec_87 : _GEN_6656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6658 = 7'h58 == _myNewVec_77_T_3[6:0] ? myVec_88 : _GEN_6657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6659 = 7'h59 == _myNewVec_77_T_3[6:0] ? myVec_89 : _GEN_6658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6660 = 7'h5a == _myNewVec_77_T_3[6:0] ? myVec_90 : _GEN_6659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6661 = 7'h5b == _myNewVec_77_T_3[6:0] ? myVec_91 : _GEN_6660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6662 = 7'h5c == _myNewVec_77_T_3[6:0] ? myVec_92 : _GEN_6661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6663 = 7'h5d == _myNewVec_77_T_3[6:0] ? myVec_93 : _GEN_6662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6664 = 7'h5e == _myNewVec_77_T_3[6:0] ? myVec_94 : _GEN_6663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6665 = 7'h5f == _myNewVec_77_T_3[6:0] ? myVec_95 : _GEN_6664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6666 = 7'h60 == _myNewVec_77_T_3[6:0] ? myVec_96 : _GEN_6665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6667 = 7'h61 == _myNewVec_77_T_3[6:0] ? myVec_97 : _GEN_6666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6668 = 7'h62 == _myNewVec_77_T_3[6:0] ? myVec_98 : _GEN_6667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6669 = 7'h63 == _myNewVec_77_T_3[6:0] ? myVec_99 : _GEN_6668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6670 = 7'h64 == _myNewVec_77_T_3[6:0] ? myVec_100 : _GEN_6669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6671 = 7'h65 == _myNewVec_77_T_3[6:0] ? myVec_101 : _GEN_6670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6672 = 7'h66 == _myNewVec_77_T_3[6:0] ? myVec_102 : _GEN_6671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6673 = 7'h67 == _myNewVec_77_T_3[6:0] ? myVec_103 : _GEN_6672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6674 = 7'h68 == _myNewVec_77_T_3[6:0] ? myVec_104 : _GEN_6673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6675 = 7'h69 == _myNewVec_77_T_3[6:0] ? myVec_105 : _GEN_6674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6676 = 7'h6a == _myNewVec_77_T_3[6:0] ? myVec_106 : _GEN_6675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6677 = 7'h6b == _myNewVec_77_T_3[6:0] ? myVec_107 : _GEN_6676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6678 = 7'h6c == _myNewVec_77_T_3[6:0] ? myVec_108 : _GEN_6677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6679 = 7'h6d == _myNewVec_77_T_3[6:0] ? myVec_109 : _GEN_6678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6680 = 7'h6e == _myNewVec_77_T_3[6:0] ? myVec_110 : _GEN_6679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6681 = 7'h6f == _myNewVec_77_T_3[6:0] ? myVec_111 : _GEN_6680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6682 = 7'h70 == _myNewVec_77_T_3[6:0] ? myVec_112 : _GEN_6681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6683 = 7'h71 == _myNewVec_77_T_3[6:0] ? myVec_113 : _GEN_6682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6684 = 7'h72 == _myNewVec_77_T_3[6:0] ? myVec_114 : _GEN_6683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6685 = 7'h73 == _myNewVec_77_T_3[6:0] ? myVec_115 : _GEN_6684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6686 = 7'h74 == _myNewVec_77_T_3[6:0] ? myVec_116 : _GEN_6685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6687 = 7'h75 == _myNewVec_77_T_3[6:0] ? myVec_117 : _GEN_6686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6688 = 7'h76 == _myNewVec_77_T_3[6:0] ? myVec_118 : _GEN_6687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6689 = 7'h77 == _myNewVec_77_T_3[6:0] ? myVec_119 : _GEN_6688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6690 = 7'h78 == _myNewVec_77_T_3[6:0] ? myVec_120 : _GEN_6689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6691 = 7'h79 == _myNewVec_77_T_3[6:0] ? myVec_121 : _GEN_6690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6692 = 7'h7a == _myNewVec_77_T_3[6:0] ? myVec_122 : _GEN_6691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6693 = 7'h7b == _myNewVec_77_T_3[6:0] ? myVec_123 : _GEN_6692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6694 = 7'h7c == _myNewVec_77_T_3[6:0] ? myVec_124 : _GEN_6693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6695 = 7'h7d == _myNewVec_77_T_3[6:0] ? myVec_125 : _GEN_6694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6696 = 7'h7e == _myNewVec_77_T_3[6:0] ? myVec_126 : _GEN_6695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_77 = 7'h7f == _myNewVec_77_T_3[6:0] ? myVec_127 : _GEN_6696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_76_T_3 = _myNewVec_127_T_1 + 16'h33; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_6699 = 7'h1 == _myNewVec_76_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6700 = 7'h2 == _myNewVec_76_T_3[6:0] ? myVec_2 : _GEN_6699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6701 = 7'h3 == _myNewVec_76_T_3[6:0] ? myVec_3 : _GEN_6700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6702 = 7'h4 == _myNewVec_76_T_3[6:0] ? myVec_4 : _GEN_6701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6703 = 7'h5 == _myNewVec_76_T_3[6:0] ? myVec_5 : _GEN_6702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6704 = 7'h6 == _myNewVec_76_T_3[6:0] ? myVec_6 : _GEN_6703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6705 = 7'h7 == _myNewVec_76_T_3[6:0] ? myVec_7 : _GEN_6704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6706 = 7'h8 == _myNewVec_76_T_3[6:0] ? myVec_8 : _GEN_6705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6707 = 7'h9 == _myNewVec_76_T_3[6:0] ? myVec_9 : _GEN_6706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6708 = 7'ha == _myNewVec_76_T_3[6:0] ? myVec_10 : _GEN_6707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6709 = 7'hb == _myNewVec_76_T_3[6:0] ? myVec_11 : _GEN_6708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6710 = 7'hc == _myNewVec_76_T_3[6:0] ? myVec_12 : _GEN_6709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6711 = 7'hd == _myNewVec_76_T_3[6:0] ? myVec_13 : _GEN_6710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6712 = 7'he == _myNewVec_76_T_3[6:0] ? myVec_14 : _GEN_6711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6713 = 7'hf == _myNewVec_76_T_3[6:0] ? myVec_15 : _GEN_6712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6714 = 7'h10 == _myNewVec_76_T_3[6:0] ? myVec_16 : _GEN_6713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6715 = 7'h11 == _myNewVec_76_T_3[6:0] ? myVec_17 : _GEN_6714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6716 = 7'h12 == _myNewVec_76_T_3[6:0] ? myVec_18 : _GEN_6715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6717 = 7'h13 == _myNewVec_76_T_3[6:0] ? myVec_19 : _GEN_6716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6718 = 7'h14 == _myNewVec_76_T_3[6:0] ? myVec_20 : _GEN_6717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6719 = 7'h15 == _myNewVec_76_T_3[6:0] ? myVec_21 : _GEN_6718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6720 = 7'h16 == _myNewVec_76_T_3[6:0] ? myVec_22 : _GEN_6719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6721 = 7'h17 == _myNewVec_76_T_3[6:0] ? myVec_23 : _GEN_6720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6722 = 7'h18 == _myNewVec_76_T_3[6:0] ? myVec_24 : _GEN_6721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6723 = 7'h19 == _myNewVec_76_T_3[6:0] ? myVec_25 : _GEN_6722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6724 = 7'h1a == _myNewVec_76_T_3[6:0] ? myVec_26 : _GEN_6723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6725 = 7'h1b == _myNewVec_76_T_3[6:0] ? myVec_27 : _GEN_6724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6726 = 7'h1c == _myNewVec_76_T_3[6:0] ? myVec_28 : _GEN_6725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6727 = 7'h1d == _myNewVec_76_T_3[6:0] ? myVec_29 : _GEN_6726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6728 = 7'h1e == _myNewVec_76_T_3[6:0] ? myVec_30 : _GEN_6727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6729 = 7'h1f == _myNewVec_76_T_3[6:0] ? myVec_31 : _GEN_6728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6730 = 7'h20 == _myNewVec_76_T_3[6:0] ? myVec_32 : _GEN_6729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6731 = 7'h21 == _myNewVec_76_T_3[6:0] ? myVec_33 : _GEN_6730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6732 = 7'h22 == _myNewVec_76_T_3[6:0] ? myVec_34 : _GEN_6731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6733 = 7'h23 == _myNewVec_76_T_3[6:0] ? myVec_35 : _GEN_6732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6734 = 7'h24 == _myNewVec_76_T_3[6:0] ? myVec_36 : _GEN_6733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6735 = 7'h25 == _myNewVec_76_T_3[6:0] ? myVec_37 : _GEN_6734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6736 = 7'h26 == _myNewVec_76_T_3[6:0] ? myVec_38 : _GEN_6735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6737 = 7'h27 == _myNewVec_76_T_3[6:0] ? myVec_39 : _GEN_6736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6738 = 7'h28 == _myNewVec_76_T_3[6:0] ? myVec_40 : _GEN_6737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6739 = 7'h29 == _myNewVec_76_T_3[6:0] ? myVec_41 : _GEN_6738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6740 = 7'h2a == _myNewVec_76_T_3[6:0] ? myVec_42 : _GEN_6739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6741 = 7'h2b == _myNewVec_76_T_3[6:0] ? myVec_43 : _GEN_6740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6742 = 7'h2c == _myNewVec_76_T_3[6:0] ? myVec_44 : _GEN_6741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6743 = 7'h2d == _myNewVec_76_T_3[6:0] ? myVec_45 : _GEN_6742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6744 = 7'h2e == _myNewVec_76_T_3[6:0] ? myVec_46 : _GEN_6743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6745 = 7'h2f == _myNewVec_76_T_3[6:0] ? myVec_47 : _GEN_6744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6746 = 7'h30 == _myNewVec_76_T_3[6:0] ? myVec_48 : _GEN_6745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6747 = 7'h31 == _myNewVec_76_T_3[6:0] ? myVec_49 : _GEN_6746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6748 = 7'h32 == _myNewVec_76_T_3[6:0] ? myVec_50 : _GEN_6747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6749 = 7'h33 == _myNewVec_76_T_3[6:0] ? myVec_51 : _GEN_6748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6750 = 7'h34 == _myNewVec_76_T_3[6:0] ? myVec_52 : _GEN_6749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6751 = 7'h35 == _myNewVec_76_T_3[6:0] ? myVec_53 : _GEN_6750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6752 = 7'h36 == _myNewVec_76_T_3[6:0] ? myVec_54 : _GEN_6751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6753 = 7'h37 == _myNewVec_76_T_3[6:0] ? myVec_55 : _GEN_6752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6754 = 7'h38 == _myNewVec_76_T_3[6:0] ? myVec_56 : _GEN_6753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6755 = 7'h39 == _myNewVec_76_T_3[6:0] ? myVec_57 : _GEN_6754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6756 = 7'h3a == _myNewVec_76_T_3[6:0] ? myVec_58 : _GEN_6755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6757 = 7'h3b == _myNewVec_76_T_3[6:0] ? myVec_59 : _GEN_6756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6758 = 7'h3c == _myNewVec_76_T_3[6:0] ? myVec_60 : _GEN_6757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6759 = 7'h3d == _myNewVec_76_T_3[6:0] ? myVec_61 : _GEN_6758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6760 = 7'h3e == _myNewVec_76_T_3[6:0] ? myVec_62 : _GEN_6759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6761 = 7'h3f == _myNewVec_76_T_3[6:0] ? myVec_63 : _GEN_6760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6762 = 7'h40 == _myNewVec_76_T_3[6:0] ? myVec_64 : _GEN_6761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6763 = 7'h41 == _myNewVec_76_T_3[6:0] ? myVec_65 : _GEN_6762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6764 = 7'h42 == _myNewVec_76_T_3[6:0] ? myVec_66 : _GEN_6763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6765 = 7'h43 == _myNewVec_76_T_3[6:0] ? myVec_67 : _GEN_6764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6766 = 7'h44 == _myNewVec_76_T_3[6:0] ? myVec_68 : _GEN_6765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6767 = 7'h45 == _myNewVec_76_T_3[6:0] ? myVec_69 : _GEN_6766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6768 = 7'h46 == _myNewVec_76_T_3[6:0] ? myVec_70 : _GEN_6767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6769 = 7'h47 == _myNewVec_76_T_3[6:0] ? myVec_71 : _GEN_6768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6770 = 7'h48 == _myNewVec_76_T_3[6:0] ? myVec_72 : _GEN_6769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6771 = 7'h49 == _myNewVec_76_T_3[6:0] ? myVec_73 : _GEN_6770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6772 = 7'h4a == _myNewVec_76_T_3[6:0] ? myVec_74 : _GEN_6771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6773 = 7'h4b == _myNewVec_76_T_3[6:0] ? myVec_75 : _GEN_6772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6774 = 7'h4c == _myNewVec_76_T_3[6:0] ? myVec_76 : _GEN_6773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6775 = 7'h4d == _myNewVec_76_T_3[6:0] ? myVec_77 : _GEN_6774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6776 = 7'h4e == _myNewVec_76_T_3[6:0] ? myVec_78 : _GEN_6775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6777 = 7'h4f == _myNewVec_76_T_3[6:0] ? myVec_79 : _GEN_6776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6778 = 7'h50 == _myNewVec_76_T_3[6:0] ? myVec_80 : _GEN_6777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6779 = 7'h51 == _myNewVec_76_T_3[6:0] ? myVec_81 : _GEN_6778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6780 = 7'h52 == _myNewVec_76_T_3[6:0] ? myVec_82 : _GEN_6779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6781 = 7'h53 == _myNewVec_76_T_3[6:0] ? myVec_83 : _GEN_6780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6782 = 7'h54 == _myNewVec_76_T_3[6:0] ? myVec_84 : _GEN_6781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6783 = 7'h55 == _myNewVec_76_T_3[6:0] ? myVec_85 : _GEN_6782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6784 = 7'h56 == _myNewVec_76_T_3[6:0] ? myVec_86 : _GEN_6783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6785 = 7'h57 == _myNewVec_76_T_3[6:0] ? myVec_87 : _GEN_6784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6786 = 7'h58 == _myNewVec_76_T_3[6:0] ? myVec_88 : _GEN_6785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6787 = 7'h59 == _myNewVec_76_T_3[6:0] ? myVec_89 : _GEN_6786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6788 = 7'h5a == _myNewVec_76_T_3[6:0] ? myVec_90 : _GEN_6787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6789 = 7'h5b == _myNewVec_76_T_3[6:0] ? myVec_91 : _GEN_6788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6790 = 7'h5c == _myNewVec_76_T_3[6:0] ? myVec_92 : _GEN_6789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6791 = 7'h5d == _myNewVec_76_T_3[6:0] ? myVec_93 : _GEN_6790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6792 = 7'h5e == _myNewVec_76_T_3[6:0] ? myVec_94 : _GEN_6791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6793 = 7'h5f == _myNewVec_76_T_3[6:0] ? myVec_95 : _GEN_6792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6794 = 7'h60 == _myNewVec_76_T_3[6:0] ? myVec_96 : _GEN_6793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6795 = 7'h61 == _myNewVec_76_T_3[6:0] ? myVec_97 : _GEN_6794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6796 = 7'h62 == _myNewVec_76_T_3[6:0] ? myVec_98 : _GEN_6795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6797 = 7'h63 == _myNewVec_76_T_3[6:0] ? myVec_99 : _GEN_6796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6798 = 7'h64 == _myNewVec_76_T_3[6:0] ? myVec_100 : _GEN_6797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6799 = 7'h65 == _myNewVec_76_T_3[6:0] ? myVec_101 : _GEN_6798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6800 = 7'h66 == _myNewVec_76_T_3[6:0] ? myVec_102 : _GEN_6799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6801 = 7'h67 == _myNewVec_76_T_3[6:0] ? myVec_103 : _GEN_6800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6802 = 7'h68 == _myNewVec_76_T_3[6:0] ? myVec_104 : _GEN_6801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6803 = 7'h69 == _myNewVec_76_T_3[6:0] ? myVec_105 : _GEN_6802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6804 = 7'h6a == _myNewVec_76_T_3[6:0] ? myVec_106 : _GEN_6803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6805 = 7'h6b == _myNewVec_76_T_3[6:0] ? myVec_107 : _GEN_6804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6806 = 7'h6c == _myNewVec_76_T_3[6:0] ? myVec_108 : _GEN_6805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6807 = 7'h6d == _myNewVec_76_T_3[6:0] ? myVec_109 : _GEN_6806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6808 = 7'h6e == _myNewVec_76_T_3[6:0] ? myVec_110 : _GEN_6807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6809 = 7'h6f == _myNewVec_76_T_3[6:0] ? myVec_111 : _GEN_6808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6810 = 7'h70 == _myNewVec_76_T_3[6:0] ? myVec_112 : _GEN_6809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6811 = 7'h71 == _myNewVec_76_T_3[6:0] ? myVec_113 : _GEN_6810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6812 = 7'h72 == _myNewVec_76_T_3[6:0] ? myVec_114 : _GEN_6811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6813 = 7'h73 == _myNewVec_76_T_3[6:0] ? myVec_115 : _GEN_6812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6814 = 7'h74 == _myNewVec_76_T_3[6:0] ? myVec_116 : _GEN_6813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6815 = 7'h75 == _myNewVec_76_T_3[6:0] ? myVec_117 : _GEN_6814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6816 = 7'h76 == _myNewVec_76_T_3[6:0] ? myVec_118 : _GEN_6815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6817 = 7'h77 == _myNewVec_76_T_3[6:0] ? myVec_119 : _GEN_6816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6818 = 7'h78 == _myNewVec_76_T_3[6:0] ? myVec_120 : _GEN_6817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6819 = 7'h79 == _myNewVec_76_T_3[6:0] ? myVec_121 : _GEN_6818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6820 = 7'h7a == _myNewVec_76_T_3[6:0] ? myVec_122 : _GEN_6819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6821 = 7'h7b == _myNewVec_76_T_3[6:0] ? myVec_123 : _GEN_6820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6822 = 7'h7c == _myNewVec_76_T_3[6:0] ? myVec_124 : _GEN_6821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6823 = 7'h7d == _myNewVec_76_T_3[6:0] ? myVec_125 : _GEN_6822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6824 = 7'h7e == _myNewVec_76_T_3[6:0] ? myVec_126 : _GEN_6823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_76 = 7'h7f == _myNewVec_76_T_3[6:0] ? myVec_127 : _GEN_6824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_75_T_3 = _myNewVec_127_T_1 + 16'h34; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_6827 = 7'h1 == _myNewVec_75_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6828 = 7'h2 == _myNewVec_75_T_3[6:0] ? myVec_2 : _GEN_6827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6829 = 7'h3 == _myNewVec_75_T_3[6:0] ? myVec_3 : _GEN_6828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6830 = 7'h4 == _myNewVec_75_T_3[6:0] ? myVec_4 : _GEN_6829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6831 = 7'h5 == _myNewVec_75_T_3[6:0] ? myVec_5 : _GEN_6830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6832 = 7'h6 == _myNewVec_75_T_3[6:0] ? myVec_6 : _GEN_6831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6833 = 7'h7 == _myNewVec_75_T_3[6:0] ? myVec_7 : _GEN_6832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6834 = 7'h8 == _myNewVec_75_T_3[6:0] ? myVec_8 : _GEN_6833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6835 = 7'h9 == _myNewVec_75_T_3[6:0] ? myVec_9 : _GEN_6834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6836 = 7'ha == _myNewVec_75_T_3[6:0] ? myVec_10 : _GEN_6835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6837 = 7'hb == _myNewVec_75_T_3[6:0] ? myVec_11 : _GEN_6836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6838 = 7'hc == _myNewVec_75_T_3[6:0] ? myVec_12 : _GEN_6837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6839 = 7'hd == _myNewVec_75_T_3[6:0] ? myVec_13 : _GEN_6838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6840 = 7'he == _myNewVec_75_T_3[6:0] ? myVec_14 : _GEN_6839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6841 = 7'hf == _myNewVec_75_T_3[6:0] ? myVec_15 : _GEN_6840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6842 = 7'h10 == _myNewVec_75_T_3[6:0] ? myVec_16 : _GEN_6841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6843 = 7'h11 == _myNewVec_75_T_3[6:0] ? myVec_17 : _GEN_6842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6844 = 7'h12 == _myNewVec_75_T_3[6:0] ? myVec_18 : _GEN_6843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6845 = 7'h13 == _myNewVec_75_T_3[6:0] ? myVec_19 : _GEN_6844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6846 = 7'h14 == _myNewVec_75_T_3[6:0] ? myVec_20 : _GEN_6845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6847 = 7'h15 == _myNewVec_75_T_3[6:0] ? myVec_21 : _GEN_6846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6848 = 7'h16 == _myNewVec_75_T_3[6:0] ? myVec_22 : _GEN_6847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6849 = 7'h17 == _myNewVec_75_T_3[6:0] ? myVec_23 : _GEN_6848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6850 = 7'h18 == _myNewVec_75_T_3[6:0] ? myVec_24 : _GEN_6849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6851 = 7'h19 == _myNewVec_75_T_3[6:0] ? myVec_25 : _GEN_6850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6852 = 7'h1a == _myNewVec_75_T_3[6:0] ? myVec_26 : _GEN_6851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6853 = 7'h1b == _myNewVec_75_T_3[6:0] ? myVec_27 : _GEN_6852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6854 = 7'h1c == _myNewVec_75_T_3[6:0] ? myVec_28 : _GEN_6853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6855 = 7'h1d == _myNewVec_75_T_3[6:0] ? myVec_29 : _GEN_6854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6856 = 7'h1e == _myNewVec_75_T_3[6:0] ? myVec_30 : _GEN_6855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6857 = 7'h1f == _myNewVec_75_T_3[6:0] ? myVec_31 : _GEN_6856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6858 = 7'h20 == _myNewVec_75_T_3[6:0] ? myVec_32 : _GEN_6857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6859 = 7'h21 == _myNewVec_75_T_3[6:0] ? myVec_33 : _GEN_6858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6860 = 7'h22 == _myNewVec_75_T_3[6:0] ? myVec_34 : _GEN_6859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6861 = 7'h23 == _myNewVec_75_T_3[6:0] ? myVec_35 : _GEN_6860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6862 = 7'h24 == _myNewVec_75_T_3[6:0] ? myVec_36 : _GEN_6861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6863 = 7'h25 == _myNewVec_75_T_3[6:0] ? myVec_37 : _GEN_6862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6864 = 7'h26 == _myNewVec_75_T_3[6:0] ? myVec_38 : _GEN_6863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6865 = 7'h27 == _myNewVec_75_T_3[6:0] ? myVec_39 : _GEN_6864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6866 = 7'h28 == _myNewVec_75_T_3[6:0] ? myVec_40 : _GEN_6865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6867 = 7'h29 == _myNewVec_75_T_3[6:0] ? myVec_41 : _GEN_6866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6868 = 7'h2a == _myNewVec_75_T_3[6:0] ? myVec_42 : _GEN_6867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6869 = 7'h2b == _myNewVec_75_T_3[6:0] ? myVec_43 : _GEN_6868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6870 = 7'h2c == _myNewVec_75_T_3[6:0] ? myVec_44 : _GEN_6869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6871 = 7'h2d == _myNewVec_75_T_3[6:0] ? myVec_45 : _GEN_6870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6872 = 7'h2e == _myNewVec_75_T_3[6:0] ? myVec_46 : _GEN_6871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6873 = 7'h2f == _myNewVec_75_T_3[6:0] ? myVec_47 : _GEN_6872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6874 = 7'h30 == _myNewVec_75_T_3[6:0] ? myVec_48 : _GEN_6873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6875 = 7'h31 == _myNewVec_75_T_3[6:0] ? myVec_49 : _GEN_6874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6876 = 7'h32 == _myNewVec_75_T_3[6:0] ? myVec_50 : _GEN_6875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6877 = 7'h33 == _myNewVec_75_T_3[6:0] ? myVec_51 : _GEN_6876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6878 = 7'h34 == _myNewVec_75_T_3[6:0] ? myVec_52 : _GEN_6877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6879 = 7'h35 == _myNewVec_75_T_3[6:0] ? myVec_53 : _GEN_6878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6880 = 7'h36 == _myNewVec_75_T_3[6:0] ? myVec_54 : _GEN_6879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6881 = 7'h37 == _myNewVec_75_T_3[6:0] ? myVec_55 : _GEN_6880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6882 = 7'h38 == _myNewVec_75_T_3[6:0] ? myVec_56 : _GEN_6881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6883 = 7'h39 == _myNewVec_75_T_3[6:0] ? myVec_57 : _GEN_6882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6884 = 7'h3a == _myNewVec_75_T_3[6:0] ? myVec_58 : _GEN_6883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6885 = 7'h3b == _myNewVec_75_T_3[6:0] ? myVec_59 : _GEN_6884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6886 = 7'h3c == _myNewVec_75_T_3[6:0] ? myVec_60 : _GEN_6885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6887 = 7'h3d == _myNewVec_75_T_3[6:0] ? myVec_61 : _GEN_6886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6888 = 7'h3e == _myNewVec_75_T_3[6:0] ? myVec_62 : _GEN_6887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6889 = 7'h3f == _myNewVec_75_T_3[6:0] ? myVec_63 : _GEN_6888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6890 = 7'h40 == _myNewVec_75_T_3[6:0] ? myVec_64 : _GEN_6889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6891 = 7'h41 == _myNewVec_75_T_3[6:0] ? myVec_65 : _GEN_6890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6892 = 7'h42 == _myNewVec_75_T_3[6:0] ? myVec_66 : _GEN_6891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6893 = 7'h43 == _myNewVec_75_T_3[6:0] ? myVec_67 : _GEN_6892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6894 = 7'h44 == _myNewVec_75_T_3[6:0] ? myVec_68 : _GEN_6893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6895 = 7'h45 == _myNewVec_75_T_3[6:0] ? myVec_69 : _GEN_6894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6896 = 7'h46 == _myNewVec_75_T_3[6:0] ? myVec_70 : _GEN_6895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6897 = 7'h47 == _myNewVec_75_T_3[6:0] ? myVec_71 : _GEN_6896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6898 = 7'h48 == _myNewVec_75_T_3[6:0] ? myVec_72 : _GEN_6897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6899 = 7'h49 == _myNewVec_75_T_3[6:0] ? myVec_73 : _GEN_6898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6900 = 7'h4a == _myNewVec_75_T_3[6:0] ? myVec_74 : _GEN_6899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6901 = 7'h4b == _myNewVec_75_T_3[6:0] ? myVec_75 : _GEN_6900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6902 = 7'h4c == _myNewVec_75_T_3[6:0] ? myVec_76 : _GEN_6901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6903 = 7'h4d == _myNewVec_75_T_3[6:0] ? myVec_77 : _GEN_6902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6904 = 7'h4e == _myNewVec_75_T_3[6:0] ? myVec_78 : _GEN_6903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6905 = 7'h4f == _myNewVec_75_T_3[6:0] ? myVec_79 : _GEN_6904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6906 = 7'h50 == _myNewVec_75_T_3[6:0] ? myVec_80 : _GEN_6905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6907 = 7'h51 == _myNewVec_75_T_3[6:0] ? myVec_81 : _GEN_6906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6908 = 7'h52 == _myNewVec_75_T_3[6:0] ? myVec_82 : _GEN_6907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6909 = 7'h53 == _myNewVec_75_T_3[6:0] ? myVec_83 : _GEN_6908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6910 = 7'h54 == _myNewVec_75_T_3[6:0] ? myVec_84 : _GEN_6909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6911 = 7'h55 == _myNewVec_75_T_3[6:0] ? myVec_85 : _GEN_6910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6912 = 7'h56 == _myNewVec_75_T_3[6:0] ? myVec_86 : _GEN_6911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6913 = 7'h57 == _myNewVec_75_T_3[6:0] ? myVec_87 : _GEN_6912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6914 = 7'h58 == _myNewVec_75_T_3[6:0] ? myVec_88 : _GEN_6913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6915 = 7'h59 == _myNewVec_75_T_3[6:0] ? myVec_89 : _GEN_6914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6916 = 7'h5a == _myNewVec_75_T_3[6:0] ? myVec_90 : _GEN_6915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6917 = 7'h5b == _myNewVec_75_T_3[6:0] ? myVec_91 : _GEN_6916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6918 = 7'h5c == _myNewVec_75_T_3[6:0] ? myVec_92 : _GEN_6917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6919 = 7'h5d == _myNewVec_75_T_3[6:0] ? myVec_93 : _GEN_6918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6920 = 7'h5e == _myNewVec_75_T_3[6:0] ? myVec_94 : _GEN_6919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6921 = 7'h5f == _myNewVec_75_T_3[6:0] ? myVec_95 : _GEN_6920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6922 = 7'h60 == _myNewVec_75_T_3[6:0] ? myVec_96 : _GEN_6921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6923 = 7'h61 == _myNewVec_75_T_3[6:0] ? myVec_97 : _GEN_6922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6924 = 7'h62 == _myNewVec_75_T_3[6:0] ? myVec_98 : _GEN_6923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6925 = 7'h63 == _myNewVec_75_T_3[6:0] ? myVec_99 : _GEN_6924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6926 = 7'h64 == _myNewVec_75_T_3[6:0] ? myVec_100 : _GEN_6925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6927 = 7'h65 == _myNewVec_75_T_3[6:0] ? myVec_101 : _GEN_6926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6928 = 7'h66 == _myNewVec_75_T_3[6:0] ? myVec_102 : _GEN_6927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6929 = 7'h67 == _myNewVec_75_T_3[6:0] ? myVec_103 : _GEN_6928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6930 = 7'h68 == _myNewVec_75_T_3[6:0] ? myVec_104 : _GEN_6929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6931 = 7'h69 == _myNewVec_75_T_3[6:0] ? myVec_105 : _GEN_6930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6932 = 7'h6a == _myNewVec_75_T_3[6:0] ? myVec_106 : _GEN_6931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6933 = 7'h6b == _myNewVec_75_T_3[6:0] ? myVec_107 : _GEN_6932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6934 = 7'h6c == _myNewVec_75_T_3[6:0] ? myVec_108 : _GEN_6933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6935 = 7'h6d == _myNewVec_75_T_3[6:0] ? myVec_109 : _GEN_6934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6936 = 7'h6e == _myNewVec_75_T_3[6:0] ? myVec_110 : _GEN_6935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6937 = 7'h6f == _myNewVec_75_T_3[6:0] ? myVec_111 : _GEN_6936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6938 = 7'h70 == _myNewVec_75_T_3[6:0] ? myVec_112 : _GEN_6937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6939 = 7'h71 == _myNewVec_75_T_3[6:0] ? myVec_113 : _GEN_6938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6940 = 7'h72 == _myNewVec_75_T_3[6:0] ? myVec_114 : _GEN_6939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6941 = 7'h73 == _myNewVec_75_T_3[6:0] ? myVec_115 : _GEN_6940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6942 = 7'h74 == _myNewVec_75_T_3[6:0] ? myVec_116 : _GEN_6941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6943 = 7'h75 == _myNewVec_75_T_3[6:0] ? myVec_117 : _GEN_6942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6944 = 7'h76 == _myNewVec_75_T_3[6:0] ? myVec_118 : _GEN_6943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6945 = 7'h77 == _myNewVec_75_T_3[6:0] ? myVec_119 : _GEN_6944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6946 = 7'h78 == _myNewVec_75_T_3[6:0] ? myVec_120 : _GEN_6945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6947 = 7'h79 == _myNewVec_75_T_3[6:0] ? myVec_121 : _GEN_6946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6948 = 7'h7a == _myNewVec_75_T_3[6:0] ? myVec_122 : _GEN_6947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6949 = 7'h7b == _myNewVec_75_T_3[6:0] ? myVec_123 : _GEN_6948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6950 = 7'h7c == _myNewVec_75_T_3[6:0] ? myVec_124 : _GEN_6949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6951 = 7'h7d == _myNewVec_75_T_3[6:0] ? myVec_125 : _GEN_6950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6952 = 7'h7e == _myNewVec_75_T_3[6:0] ? myVec_126 : _GEN_6951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_75 = 7'h7f == _myNewVec_75_T_3[6:0] ? myVec_127 : _GEN_6952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_74_T_3 = _myNewVec_127_T_1 + 16'h35; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_6955 = 7'h1 == _myNewVec_74_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6956 = 7'h2 == _myNewVec_74_T_3[6:0] ? myVec_2 : _GEN_6955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6957 = 7'h3 == _myNewVec_74_T_3[6:0] ? myVec_3 : _GEN_6956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6958 = 7'h4 == _myNewVec_74_T_3[6:0] ? myVec_4 : _GEN_6957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6959 = 7'h5 == _myNewVec_74_T_3[6:0] ? myVec_5 : _GEN_6958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6960 = 7'h6 == _myNewVec_74_T_3[6:0] ? myVec_6 : _GEN_6959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6961 = 7'h7 == _myNewVec_74_T_3[6:0] ? myVec_7 : _GEN_6960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6962 = 7'h8 == _myNewVec_74_T_3[6:0] ? myVec_8 : _GEN_6961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6963 = 7'h9 == _myNewVec_74_T_3[6:0] ? myVec_9 : _GEN_6962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6964 = 7'ha == _myNewVec_74_T_3[6:0] ? myVec_10 : _GEN_6963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6965 = 7'hb == _myNewVec_74_T_3[6:0] ? myVec_11 : _GEN_6964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6966 = 7'hc == _myNewVec_74_T_3[6:0] ? myVec_12 : _GEN_6965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6967 = 7'hd == _myNewVec_74_T_3[6:0] ? myVec_13 : _GEN_6966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6968 = 7'he == _myNewVec_74_T_3[6:0] ? myVec_14 : _GEN_6967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6969 = 7'hf == _myNewVec_74_T_3[6:0] ? myVec_15 : _GEN_6968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6970 = 7'h10 == _myNewVec_74_T_3[6:0] ? myVec_16 : _GEN_6969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6971 = 7'h11 == _myNewVec_74_T_3[6:0] ? myVec_17 : _GEN_6970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6972 = 7'h12 == _myNewVec_74_T_3[6:0] ? myVec_18 : _GEN_6971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6973 = 7'h13 == _myNewVec_74_T_3[6:0] ? myVec_19 : _GEN_6972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6974 = 7'h14 == _myNewVec_74_T_3[6:0] ? myVec_20 : _GEN_6973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6975 = 7'h15 == _myNewVec_74_T_3[6:0] ? myVec_21 : _GEN_6974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6976 = 7'h16 == _myNewVec_74_T_3[6:0] ? myVec_22 : _GEN_6975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6977 = 7'h17 == _myNewVec_74_T_3[6:0] ? myVec_23 : _GEN_6976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6978 = 7'h18 == _myNewVec_74_T_3[6:0] ? myVec_24 : _GEN_6977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6979 = 7'h19 == _myNewVec_74_T_3[6:0] ? myVec_25 : _GEN_6978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6980 = 7'h1a == _myNewVec_74_T_3[6:0] ? myVec_26 : _GEN_6979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6981 = 7'h1b == _myNewVec_74_T_3[6:0] ? myVec_27 : _GEN_6980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6982 = 7'h1c == _myNewVec_74_T_3[6:0] ? myVec_28 : _GEN_6981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6983 = 7'h1d == _myNewVec_74_T_3[6:0] ? myVec_29 : _GEN_6982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6984 = 7'h1e == _myNewVec_74_T_3[6:0] ? myVec_30 : _GEN_6983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6985 = 7'h1f == _myNewVec_74_T_3[6:0] ? myVec_31 : _GEN_6984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6986 = 7'h20 == _myNewVec_74_T_3[6:0] ? myVec_32 : _GEN_6985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6987 = 7'h21 == _myNewVec_74_T_3[6:0] ? myVec_33 : _GEN_6986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6988 = 7'h22 == _myNewVec_74_T_3[6:0] ? myVec_34 : _GEN_6987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6989 = 7'h23 == _myNewVec_74_T_3[6:0] ? myVec_35 : _GEN_6988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6990 = 7'h24 == _myNewVec_74_T_3[6:0] ? myVec_36 : _GEN_6989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6991 = 7'h25 == _myNewVec_74_T_3[6:0] ? myVec_37 : _GEN_6990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6992 = 7'h26 == _myNewVec_74_T_3[6:0] ? myVec_38 : _GEN_6991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6993 = 7'h27 == _myNewVec_74_T_3[6:0] ? myVec_39 : _GEN_6992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6994 = 7'h28 == _myNewVec_74_T_3[6:0] ? myVec_40 : _GEN_6993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6995 = 7'h29 == _myNewVec_74_T_3[6:0] ? myVec_41 : _GEN_6994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6996 = 7'h2a == _myNewVec_74_T_3[6:0] ? myVec_42 : _GEN_6995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6997 = 7'h2b == _myNewVec_74_T_3[6:0] ? myVec_43 : _GEN_6996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6998 = 7'h2c == _myNewVec_74_T_3[6:0] ? myVec_44 : _GEN_6997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_6999 = 7'h2d == _myNewVec_74_T_3[6:0] ? myVec_45 : _GEN_6998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7000 = 7'h2e == _myNewVec_74_T_3[6:0] ? myVec_46 : _GEN_6999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7001 = 7'h2f == _myNewVec_74_T_3[6:0] ? myVec_47 : _GEN_7000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7002 = 7'h30 == _myNewVec_74_T_3[6:0] ? myVec_48 : _GEN_7001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7003 = 7'h31 == _myNewVec_74_T_3[6:0] ? myVec_49 : _GEN_7002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7004 = 7'h32 == _myNewVec_74_T_3[6:0] ? myVec_50 : _GEN_7003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7005 = 7'h33 == _myNewVec_74_T_3[6:0] ? myVec_51 : _GEN_7004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7006 = 7'h34 == _myNewVec_74_T_3[6:0] ? myVec_52 : _GEN_7005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7007 = 7'h35 == _myNewVec_74_T_3[6:0] ? myVec_53 : _GEN_7006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7008 = 7'h36 == _myNewVec_74_T_3[6:0] ? myVec_54 : _GEN_7007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7009 = 7'h37 == _myNewVec_74_T_3[6:0] ? myVec_55 : _GEN_7008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7010 = 7'h38 == _myNewVec_74_T_3[6:0] ? myVec_56 : _GEN_7009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7011 = 7'h39 == _myNewVec_74_T_3[6:0] ? myVec_57 : _GEN_7010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7012 = 7'h3a == _myNewVec_74_T_3[6:0] ? myVec_58 : _GEN_7011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7013 = 7'h3b == _myNewVec_74_T_3[6:0] ? myVec_59 : _GEN_7012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7014 = 7'h3c == _myNewVec_74_T_3[6:0] ? myVec_60 : _GEN_7013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7015 = 7'h3d == _myNewVec_74_T_3[6:0] ? myVec_61 : _GEN_7014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7016 = 7'h3e == _myNewVec_74_T_3[6:0] ? myVec_62 : _GEN_7015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7017 = 7'h3f == _myNewVec_74_T_3[6:0] ? myVec_63 : _GEN_7016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7018 = 7'h40 == _myNewVec_74_T_3[6:0] ? myVec_64 : _GEN_7017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7019 = 7'h41 == _myNewVec_74_T_3[6:0] ? myVec_65 : _GEN_7018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7020 = 7'h42 == _myNewVec_74_T_3[6:0] ? myVec_66 : _GEN_7019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7021 = 7'h43 == _myNewVec_74_T_3[6:0] ? myVec_67 : _GEN_7020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7022 = 7'h44 == _myNewVec_74_T_3[6:0] ? myVec_68 : _GEN_7021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7023 = 7'h45 == _myNewVec_74_T_3[6:0] ? myVec_69 : _GEN_7022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7024 = 7'h46 == _myNewVec_74_T_3[6:0] ? myVec_70 : _GEN_7023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7025 = 7'h47 == _myNewVec_74_T_3[6:0] ? myVec_71 : _GEN_7024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7026 = 7'h48 == _myNewVec_74_T_3[6:0] ? myVec_72 : _GEN_7025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7027 = 7'h49 == _myNewVec_74_T_3[6:0] ? myVec_73 : _GEN_7026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7028 = 7'h4a == _myNewVec_74_T_3[6:0] ? myVec_74 : _GEN_7027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7029 = 7'h4b == _myNewVec_74_T_3[6:0] ? myVec_75 : _GEN_7028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7030 = 7'h4c == _myNewVec_74_T_3[6:0] ? myVec_76 : _GEN_7029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7031 = 7'h4d == _myNewVec_74_T_3[6:0] ? myVec_77 : _GEN_7030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7032 = 7'h4e == _myNewVec_74_T_3[6:0] ? myVec_78 : _GEN_7031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7033 = 7'h4f == _myNewVec_74_T_3[6:0] ? myVec_79 : _GEN_7032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7034 = 7'h50 == _myNewVec_74_T_3[6:0] ? myVec_80 : _GEN_7033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7035 = 7'h51 == _myNewVec_74_T_3[6:0] ? myVec_81 : _GEN_7034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7036 = 7'h52 == _myNewVec_74_T_3[6:0] ? myVec_82 : _GEN_7035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7037 = 7'h53 == _myNewVec_74_T_3[6:0] ? myVec_83 : _GEN_7036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7038 = 7'h54 == _myNewVec_74_T_3[6:0] ? myVec_84 : _GEN_7037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7039 = 7'h55 == _myNewVec_74_T_3[6:0] ? myVec_85 : _GEN_7038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7040 = 7'h56 == _myNewVec_74_T_3[6:0] ? myVec_86 : _GEN_7039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7041 = 7'h57 == _myNewVec_74_T_3[6:0] ? myVec_87 : _GEN_7040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7042 = 7'h58 == _myNewVec_74_T_3[6:0] ? myVec_88 : _GEN_7041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7043 = 7'h59 == _myNewVec_74_T_3[6:0] ? myVec_89 : _GEN_7042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7044 = 7'h5a == _myNewVec_74_T_3[6:0] ? myVec_90 : _GEN_7043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7045 = 7'h5b == _myNewVec_74_T_3[6:0] ? myVec_91 : _GEN_7044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7046 = 7'h5c == _myNewVec_74_T_3[6:0] ? myVec_92 : _GEN_7045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7047 = 7'h5d == _myNewVec_74_T_3[6:0] ? myVec_93 : _GEN_7046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7048 = 7'h5e == _myNewVec_74_T_3[6:0] ? myVec_94 : _GEN_7047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7049 = 7'h5f == _myNewVec_74_T_3[6:0] ? myVec_95 : _GEN_7048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7050 = 7'h60 == _myNewVec_74_T_3[6:0] ? myVec_96 : _GEN_7049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7051 = 7'h61 == _myNewVec_74_T_3[6:0] ? myVec_97 : _GEN_7050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7052 = 7'h62 == _myNewVec_74_T_3[6:0] ? myVec_98 : _GEN_7051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7053 = 7'h63 == _myNewVec_74_T_3[6:0] ? myVec_99 : _GEN_7052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7054 = 7'h64 == _myNewVec_74_T_3[6:0] ? myVec_100 : _GEN_7053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7055 = 7'h65 == _myNewVec_74_T_3[6:0] ? myVec_101 : _GEN_7054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7056 = 7'h66 == _myNewVec_74_T_3[6:0] ? myVec_102 : _GEN_7055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7057 = 7'h67 == _myNewVec_74_T_3[6:0] ? myVec_103 : _GEN_7056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7058 = 7'h68 == _myNewVec_74_T_3[6:0] ? myVec_104 : _GEN_7057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7059 = 7'h69 == _myNewVec_74_T_3[6:0] ? myVec_105 : _GEN_7058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7060 = 7'h6a == _myNewVec_74_T_3[6:0] ? myVec_106 : _GEN_7059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7061 = 7'h6b == _myNewVec_74_T_3[6:0] ? myVec_107 : _GEN_7060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7062 = 7'h6c == _myNewVec_74_T_3[6:0] ? myVec_108 : _GEN_7061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7063 = 7'h6d == _myNewVec_74_T_3[6:0] ? myVec_109 : _GEN_7062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7064 = 7'h6e == _myNewVec_74_T_3[6:0] ? myVec_110 : _GEN_7063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7065 = 7'h6f == _myNewVec_74_T_3[6:0] ? myVec_111 : _GEN_7064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7066 = 7'h70 == _myNewVec_74_T_3[6:0] ? myVec_112 : _GEN_7065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7067 = 7'h71 == _myNewVec_74_T_3[6:0] ? myVec_113 : _GEN_7066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7068 = 7'h72 == _myNewVec_74_T_3[6:0] ? myVec_114 : _GEN_7067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7069 = 7'h73 == _myNewVec_74_T_3[6:0] ? myVec_115 : _GEN_7068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7070 = 7'h74 == _myNewVec_74_T_3[6:0] ? myVec_116 : _GEN_7069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7071 = 7'h75 == _myNewVec_74_T_3[6:0] ? myVec_117 : _GEN_7070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7072 = 7'h76 == _myNewVec_74_T_3[6:0] ? myVec_118 : _GEN_7071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7073 = 7'h77 == _myNewVec_74_T_3[6:0] ? myVec_119 : _GEN_7072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7074 = 7'h78 == _myNewVec_74_T_3[6:0] ? myVec_120 : _GEN_7073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7075 = 7'h79 == _myNewVec_74_T_3[6:0] ? myVec_121 : _GEN_7074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7076 = 7'h7a == _myNewVec_74_T_3[6:0] ? myVec_122 : _GEN_7075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7077 = 7'h7b == _myNewVec_74_T_3[6:0] ? myVec_123 : _GEN_7076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7078 = 7'h7c == _myNewVec_74_T_3[6:0] ? myVec_124 : _GEN_7077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7079 = 7'h7d == _myNewVec_74_T_3[6:0] ? myVec_125 : _GEN_7078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7080 = 7'h7e == _myNewVec_74_T_3[6:0] ? myVec_126 : _GEN_7079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_74 = 7'h7f == _myNewVec_74_T_3[6:0] ? myVec_127 : _GEN_7080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_73_T_3 = _myNewVec_127_T_1 + 16'h36; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_7083 = 7'h1 == _myNewVec_73_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7084 = 7'h2 == _myNewVec_73_T_3[6:0] ? myVec_2 : _GEN_7083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7085 = 7'h3 == _myNewVec_73_T_3[6:0] ? myVec_3 : _GEN_7084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7086 = 7'h4 == _myNewVec_73_T_3[6:0] ? myVec_4 : _GEN_7085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7087 = 7'h5 == _myNewVec_73_T_3[6:0] ? myVec_5 : _GEN_7086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7088 = 7'h6 == _myNewVec_73_T_3[6:0] ? myVec_6 : _GEN_7087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7089 = 7'h7 == _myNewVec_73_T_3[6:0] ? myVec_7 : _GEN_7088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7090 = 7'h8 == _myNewVec_73_T_3[6:0] ? myVec_8 : _GEN_7089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7091 = 7'h9 == _myNewVec_73_T_3[6:0] ? myVec_9 : _GEN_7090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7092 = 7'ha == _myNewVec_73_T_3[6:0] ? myVec_10 : _GEN_7091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7093 = 7'hb == _myNewVec_73_T_3[6:0] ? myVec_11 : _GEN_7092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7094 = 7'hc == _myNewVec_73_T_3[6:0] ? myVec_12 : _GEN_7093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7095 = 7'hd == _myNewVec_73_T_3[6:0] ? myVec_13 : _GEN_7094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7096 = 7'he == _myNewVec_73_T_3[6:0] ? myVec_14 : _GEN_7095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7097 = 7'hf == _myNewVec_73_T_3[6:0] ? myVec_15 : _GEN_7096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7098 = 7'h10 == _myNewVec_73_T_3[6:0] ? myVec_16 : _GEN_7097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7099 = 7'h11 == _myNewVec_73_T_3[6:0] ? myVec_17 : _GEN_7098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7100 = 7'h12 == _myNewVec_73_T_3[6:0] ? myVec_18 : _GEN_7099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7101 = 7'h13 == _myNewVec_73_T_3[6:0] ? myVec_19 : _GEN_7100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7102 = 7'h14 == _myNewVec_73_T_3[6:0] ? myVec_20 : _GEN_7101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7103 = 7'h15 == _myNewVec_73_T_3[6:0] ? myVec_21 : _GEN_7102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7104 = 7'h16 == _myNewVec_73_T_3[6:0] ? myVec_22 : _GEN_7103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7105 = 7'h17 == _myNewVec_73_T_3[6:0] ? myVec_23 : _GEN_7104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7106 = 7'h18 == _myNewVec_73_T_3[6:0] ? myVec_24 : _GEN_7105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7107 = 7'h19 == _myNewVec_73_T_3[6:0] ? myVec_25 : _GEN_7106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7108 = 7'h1a == _myNewVec_73_T_3[6:0] ? myVec_26 : _GEN_7107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7109 = 7'h1b == _myNewVec_73_T_3[6:0] ? myVec_27 : _GEN_7108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7110 = 7'h1c == _myNewVec_73_T_3[6:0] ? myVec_28 : _GEN_7109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7111 = 7'h1d == _myNewVec_73_T_3[6:0] ? myVec_29 : _GEN_7110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7112 = 7'h1e == _myNewVec_73_T_3[6:0] ? myVec_30 : _GEN_7111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7113 = 7'h1f == _myNewVec_73_T_3[6:0] ? myVec_31 : _GEN_7112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7114 = 7'h20 == _myNewVec_73_T_3[6:0] ? myVec_32 : _GEN_7113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7115 = 7'h21 == _myNewVec_73_T_3[6:0] ? myVec_33 : _GEN_7114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7116 = 7'h22 == _myNewVec_73_T_3[6:0] ? myVec_34 : _GEN_7115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7117 = 7'h23 == _myNewVec_73_T_3[6:0] ? myVec_35 : _GEN_7116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7118 = 7'h24 == _myNewVec_73_T_3[6:0] ? myVec_36 : _GEN_7117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7119 = 7'h25 == _myNewVec_73_T_3[6:0] ? myVec_37 : _GEN_7118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7120 = 7'h26 == _myNewVec_73_T_3[6:0] ? myVec_38 : _GEN_7119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7121 = 7'h27 == _myNewVec_73_T_3[6:0] ? myVec_39 : _GEN_7120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7122 = 7'h28 == _myNewVec_73_T_3[6:0] ? myVec_40 : _GEN_7121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7123 = 7'h29 == _myNewVec_73_T_3[6:0] ? myVec_41 : _GEN_7122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7124 = 7'h2a == _myNewVec_73_T_3[6:0] ? myVec_42 : _GEN_7123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7125 = 7'h2b == _myNewVec_73_T_3[6:0] ? myVec_43 : _GEN_7124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7126 = 7'h2c == _myNewVec_73_T_3[6:0] ? myVec_44 : _GEN_7125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7127 = 7'h2d == _myNewVec_73_T_3[6:0] ? myVec_45 : _GEN_7126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7128 = 7'h2e == _myNewVec_73_T_3[6:0] ? myVec_46 : _GEN_7127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7129 = 7'h2f == _myNewVec_73_T_3[6:0] ? myVec_47 : _GEN_7128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7130 = 7'h30 == _myNewVec_73_T_3[6:0] ? myVec_48 : _GEN_7129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7131 = 7'h31 == _myNewVec_73_T_3[6:0] ? myVec_49 : _GEN_7130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7132 = 7'h32 == _myNewVec_73_T_3[6:0] ? myVec_50 : _GEN_7131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7133 = 7'h33 == _myNewVec_73_T_3[6:0] ? myVec_51 : _GEN_7132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7134 = 7'h34 == _myNewVec_73_T_3[6:0] ? myVec_52 : _GEN_7133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7135 = 7'h35 == _myNewVec_73_T_3[6:0] ? myVec_53 : _GEN_7134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7136 = 7'h36 == _myNewVec_73_T_3[6:0] ? myVec_54 : _GEN_7135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7137 = 7'h37 == _myNewVec_73_T_3[6:0] ? myVec_55 : _GEN_7136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7138 = 7'h38 == _myNewVec_73_T_3[6:0] ? myVec_56 : _GEN_7137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7139 = 7'h39 == _myNewVec_73_T_3[6:0] ? myVec_57 : _GEN_7138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7140 = 7'h3a == _myNewVec_73_T_3[6:0] ? myVec_58 : _GEN_7139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7141 = 7'h3b == _myNewVec_73_T_3[6:0] ? myVec_59 : _GEN_7140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7142 = 7'h3c == _myNewVec_73_T_3[6:0] ? myVec_60 : _GEN_7141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7143 = 7'h3d == _myNewVec_73_T_3[6:0] ? myVec_61 : _GEN_7142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7144 = 7'h3e == _myNewVec_73_T_3[6:0] ? myVec_62 : _GEN_7143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7145 = 7'h3f == _myNewVec_73_T_3[6:0] ? myVec_63 : _GEN_7144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7146 = 7'h40 == _myNewVec_73_T_3[6:0] ? myVec_64 : _GEN_7145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7147 = 7'h41 == _myNewVec_73_T_3[6:0] ? myVec_65 : _GEN_7146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7148 = 7'h42 == _myNewVec_73_T_3[6:0] ? myVec_66 : _GEN_7147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7149 = 7'h43 == _myNewVec_73_T_3[6:0] ? myVec_67 : _GEN_7148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7150 = 7'h44 == _myNewVec_73_T_3[6:0] ? myVec_68 : _GEN_7149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7151 = 7'h45 == _myNewVec_73_T_3[6:0] ? myVec_69 : _GEN_7150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7152 = 7'h46 == _myNewVec_73_T_3[6:0] ? myVec_70 : _GEN_7151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7153 = 7'h47 == _myNewVec_73_T_3[6:0] ? myVec_71 : _GEN_7152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7154 = 7'h48 == _myNewVec_73_T_3[6:0] ? myVec_72 : _GEN_7153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7155 = 7'h49 == _myNewVec_73_T_3[6:0] ? myVec_73 : _GEN_7154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7156 = 7'h4a == _myNewVec_73_T_3[6:0] ? myVec_74 : _GEN_7155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7157 = 7'h4b == _myNewVec_73_T_3[6:0] ? myVec_75 : _GEN_7156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7158 = 7'h4c == _myNewVec_73_T_3[6:0] ? myVec_76 : _GEN_7157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7159 = 7'h4d == _myNewVec_73_T_3[6:0] ? myVec_77 : _GEN_7158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7160 = 7'h4e == _myNewVec_73_T_3[6:0] ? myVec_78 : _GEN_7159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7161 = 7'h4f == _myNewVec_73_T_3[6:0] ? myVec_79 : _GEN_7160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7162 = 7'h50 == _myNewVec_73_T_3[6:0] ? myVec_80 : _GEN_7161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7163 = 7'h51 == _myNewVec_73_T_3[6:0] ? myVec_81 : _GEN_7162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7164 = 7'h52 == _myNewVec_73_T_3[6:0] ? myVec_82 : _GEN_7163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7165 = 7'h53 == _myNewVec_73_T_3[6:0] ? myVec_83 : _GEN_7164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7166 = 7'h54 == _myNewVec_73_T_3[6:0] ? myVec_84 : _GEN_7165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7167 = 7'h55 == _myNewVec_73_T_3[6:0] ? myVec_85 : _GEN_7166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7168 = 7'h56 == _myNewVec_73_T_3[6:0] ? myVec_86 : _GEN_7167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7169 = 7'h57 == _myNewVec_73_T_3[6:0] ? myVec_87 : _GEN_7168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7170 = 7'h58 == _myNewVec_73_T_3[6:0] ? myVec_88 : _GEN_7169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7171 = 7'h59 == _myNewVec_73_T_3[6:0] ? myVec_89 : _GEN_7170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7172 = 7'h5a == _myNewVec_73_T_3[6:0] ? myVec_90 : _GEN_7171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7173 = 7'h5b == _myNewVec_73_T_3[6:0] ? myVec_91 : _GEN_7172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7174 = 7'h5c == _myNewVec_73_T_3[6:0] ? myVec_92 : _GEN_7173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7175 = 7'h5d == _myNewVec_73_T_3[6:0] ? myVec_93 : _GEN_7174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7176 = 7'h5e == _myNewVec_73_T_3[6:0] ? myVec_94 : _GEN_7175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7177 = 7'h5f == _myNewVec_73_T_3[6:0] ? myVec_95 : _GEN_7176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7178 = 7'h60 == _myNewVec_73_T_3[6:0] ? myVec_96 : _GEN_7177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7179 = 7'h61 == _myNewVec_73_T_3[6:0] ? myVec_97 : _GEN_7178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7180 = 7'h62 == _myNewVec_73_T_3[6:0] ? myVec_98 : _GEN_7179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7181 = 7'h63 == _myNewVec_73_T_3[6:0] ? myVec_99 : _GEN_7180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7182 = 7'h64 == _myNewVec_73_T_3[6:0] ? myVec_100 : _GEN_7181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7183 = 7'h65 == _myNewVec_73_T_3[6:0] ? myVec_101 : _GEN_7182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7184 = 7'h66 == _myNewVec_73_T_3[6:0] ? myVec_102 : _GEN_7183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7185 = 7'h67 == _myNewVec_73_T_3[6:0] ? myVec_103 : _GEN_7184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7186 = 7'h68 == _myNewVec_73_T_3[6:0] ? myVec_104 : _GEN_7185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7187 = 7'h69 == _myNewVec_73_T_3[6:0] ? myVec_105 : _GEN_7186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7188 = 7'h6a == _myNewVec_73_T_3[6:0] ? myVec_106 : _GEN_7187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7189 = 7'h6b == _myNewVec_73_T_3[6:0] ? myVec_107 : _GEN_7188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7190 = 7'h6c == _myNewVec_73_T_3[6:0] ? myVec_108 : _GEN_7189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7191 = 7'h6d == _myNewVec_73_T_3[6:0] ? myVec_109 : _GEN_7190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7192 = 7'h6e == _myNewVec_73_T_3[6:0] ? myVec_110 : _GEN_7191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7193 = 7'h6f == _myNewVec_73_T_3[6:0] ? myVec_111 : _GEN_7192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7194 = 7'h70 == _myNewVec_73_T_3[6:0] ? myVec_112 : _GEN_7193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7195 = 7'h71 == _myNewVec_73_T_3[6:0] ? myVec_113 : _GEN_7194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7196 = 7'h72 == _myNewVec_73_T_3[6:0] ? myVec_114 : _GEN_7195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7197 = 7'h73 == _myNewVec_73_T_3[6:0] ? myVec_115 : _GEN_7196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7198 = 7'h74 == _myNewVec_73_T_3[6:0] ? myVec_116 : _GEN_7197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7199 = 7'h75 == _myNewVec_73_T_3[6:0] ? myVec_117 : _GEN_7198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7200 = 7'h76 == _myNewVec_73_T_3[6:0] ? myVec_118 : _GEN_7199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7201 = 7'h77 == _myNewVec_73_T_3[6:0] ? myVec_119 : _GEN_7200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7202 = 7'h78 == _myNewVec_73_T_3[6:0] ? myVec_120 : _GEN_7201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7203 = 7'h79 == _myNewVec_73_T_3[6:0] ? myVec_121 : _GEN_7202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7204 = 7'h7a == _myNewVec_73_T_3[6:0] ? myVec_122 : _GEN_7203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7205 = 7'h7b == _myNewVec_73_T_3[6:0] ? myVec_123 : _GEN_7204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7206 = 7'h7c == _myNewVec_73_T_3[6:0] ? myVec_124 : _GEN_7205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7207 = 7'h7d == _myNewVec_73_T_3[6:0] ? myVec_125 : _GEN_7206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7208 = 7'h7e == _myNewVec_73_T_3[6:0] ? myVec_126 : _GEN_7207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_73 = 7'h7f == _myNewVec_73_T_3[6:0] ? myVec_127 : _GEN_7208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_72_T_3 = _myNewVec_127_T_1 + 16'h37; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_7211 = 7'h1 == _myNewVec_72_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7212 = 7'h2 == _myNewVec_72_T_3[6:0] ? myVec_2 : _GEN_7211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7213 = 7'h3 == _myNewVec_72_T_3[6:0] ? myVec_3 : _GEN_7212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7214 = 7'h4 == _myNewVec_72_T_3[6:0] ? myVec_4 : _GEN_7213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7215 = 7'h5 == _myNewVec_72_T_3[6:0] ? myVec_5 : _GEN_7214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7216 = 7'h6 == _myNewVec_72_T_3[6:0] ? myVec_6 : _GEN_7215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7217 = 7'h7 == _myNewVec_72_T_3[6:0] ? myVec_7 : _GEN_7216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7218 = 7'h8 == _myNewVec_72_T_3[6:0] ? myVec_8 : _GEN_7217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7219 = 7'h9 == _myNewVec_72_T_3[6:0] ? myVec_9 : _GEN_7218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7220 = 7'ha == _myNewVec_72_T_3[6:0] ? myVec_10 : _GEN_7219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7221 = 7'hb == _myNewVec_72_T_3[6:0] ? myVec_11 : _GEN_7220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7222 = 7'hc == _myNewVec_72_T_3[6:0] ? myVec_12 : _GEN_7221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7223 = 7'hd == _myNewVec_72_T_3[6:0] ? myVec_13 : _GEN_7222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7224 = 7'he == _myNewVec_72_T_3[6:0] ? myVec_14 : _GEN_7223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7225 = 7'hf == _myNewVec_72_T_3[6:0] ? myVec_15 : _GEN_7224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7226 = 7'h10 == _myNewVec_72_T_3[6:0] ? myVec_16 : _GEN_7225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7227 = 7'h11 == _myNewVec_72_T_3[6:0] ? myVec_17 : _GEN_7226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7228 = 7'h12 == _myNewVec_72_T_3[6:0] ? myVec_18 : _GEN_7227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7229 = 7'h13 == _myNewVec_72_T_3[6:0] ? myVec_19 : _GEN_7228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7230 = 7'h14 == _myNewVec_72_T_3[6:0] ? myVec_20 : _GEN_7229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7231 = 7'h15 == _myNewVec_72_T_3[6:0] ? myVec_21 : _GEN_7230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7232 = 7'h16 == _myNewVec_72_T_3[6:0] ? myVec_22 : _GEN_7231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7233 = 7'h17 == _myNewVec_72_T_3[6:0] ? myVec_23 : _GEN_7232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7234 = 7'h18 == _myNewVec_72_T_3[6:0] ? myVec_24 : _GEN_7233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7235 = 7'h19 == _myNewVec_72_T_3[6:0] ? myVec_25 : _GEN_7234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7236 = 7'h1a == _myNewVec_72_T_3[6:0] ? myVec_26 : _GEN_7235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7237 = 7'h1b == _myNewVec_72_T_3[6:0] ? myVec_27 : _GEN_7236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7238 = 7'h1c == _myNewVec_72_T_3[6:0] ? myVec_28 : _GEN_7237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7239 = 7'h1d == _myNewVec_72_T_3[6:0] ? myVec_29 : _GEN_7238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7240 = 7'h1e == _myNewVec_72_T_3[6:0] ? myVec_30 : _GEN_7239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7241 = 7'h1f == _myNewVec_72_T_3[6:0] ? myVec_31 : _GEN_7240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7242 = 7'h20 == _myNewVec_72_T_3[6:0] ? myVec_32 : _GEN_7241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7243 = 7'h21 == _myNewVec_72_T_3[6:0] ? myVec_33 : _GEN_7242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7244 = 7'h22 == _myNewVec_72_T_3[6:0] ? myVec_34 : _GEN_7243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7245 = 7'h23 == _myNewVec_72_T_3[6:0] ? myVec_35 : _GEN_7244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7246 = 7'h24 == _myNewVec_72_T_3[6:0] ? myVec_36 : _GEN_7245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7247 = 7'h25 == _myNewVec_72_T_3[6:0] ? myVec_37 : _GEN_7246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7248 = 7'h26 == _myNewVec_72_T_3[6:0] ? myVec_38 : _GEN_7247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7249 = 7'h27 == _myNewVec_72_T_3[6:0] ? myVec_39 : _GEN_7248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7250 = 7'h28 == _myNewVec_72_T_3[6:0] ? myVec_40 : _GEN_7249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7251 = 7'h29 == _myNewVec_72_T_3[6:0] ? myVec_41 : _GEN_7250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7252 = 7'h2a == _myNewVec_72_T_3[6:0] ? myVec_42 : _GEN_7251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7253 = 7'h2b == _myNewVec_72_T_3[6:0] ? myVec_43 : _GEN_7252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7254 = 7'h2c == _myNewVec_72_T_3[6:0] ? myVec_44 : _GEN_7253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7255 = 7'h2d == _myNewVec_72_T_3[6:0] ? myVec_45 : _GEN_7254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7256 = 7'h2e == _myNewVec_72_T_3[6:0] ? myVec_46 : _GEN_7255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7257 = 7'h2f == _myNewVec_72_T_3[6:0] ? myVec_47 : _GEN_7256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7258 = 7'h30 == _myNewVec_72_T_3[6:0] ? myVec_48 : _GEN_7257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7259 = 7'h31 == _myNewVec_72_T_3[6:0] ? myVec_49 : _GEN_7258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7260 = 7'h32 == _myNewVec_72_T_3[6:0] ? myVec_50 : _GEN_7259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7261 = 7'h33 == _myNewVec_72_T_3[6:0] ? myVec_51 : _GEN_7260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7262 = 7'h34 == _myNewVec_72_T_3[6:0] ? myVec_52 : _GEN_7261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7263 = 7'h35 == _myNewVec_72_T_3[6:0] ? myVec_53 : _GEN_7262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7264 = 7'h36 == _myNewVec_72_T_3[6:0] ? myVec_54 : _GEN_7263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7265 = 7'h37 == _myNewVec_72_T_3[6:0] ? myVec_55 : _GEN_7264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7266 = 7'h38 == _myNewVec_72_T_3[6:0] ? myVec_56 : _GEN_7265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7267 = 7'h39 == _myNewVec_72_T_3[6:0] ? myVec_57 : _GEN_7266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7268 = 7'h3a == _myNewVec_72_T_3[6:0] ? myVec_58 : _GEN_7267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7269 = 7'h3b == _myNewVec_72_T_3[6:0] ? myVec_59 : _GEN_7268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7270 = 7'h3c == _myNewVec_72_T_3[6:0] ? myVec_60 : _GEN_7269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7271 = 7'h3d == _myNewVec_72_T_3[6:0] ? myVec_61 : _GEN_7270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7272 = 7'h3e == _myNewVec_72_T_3[6:0] ? myVec_62 : _GEN_7271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7273 = 7'h3f == _myNewVec_72_T_3[6:0] ? myVec_63 : _GEN_7272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7274 = 7'h40 == _myNewVec_72_T_3[6:0] ? myVec_64 : _GEN_7273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7275 = 7'h41 == _myNewVec_72_T_3[6:0] ? myVec_65 : _GEN_7274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7276 = 7'h42 == _myNewVec_72_T_3[6:0] ? myVec_66 : _GEN_7275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7277 = 7'h43 == _myNewVec_72_T_3[6:0] ? myVec_67 : _GEN_7276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7278 = 7'h44 == _myNewVec_72_T_3[6:0] ? myVec_68 : _GEN_7277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7279 = 7'h45 == _myNewVec_72_T_3[6:0] ? myVec_69 : _GEN_7278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7280 = 7'h46 == _myNewVec_72_T_3[6:0] ? myVec_70 : _GEN_7279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7281 = 7'h47 == _myNewVec_72_T_3[6:0] ? myVec_71 : _GEN_7280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7282 = 7'h48 == _myNewVec_72_T_3[6:0] ? myVec_72 : _GEN_7281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7283 = 7'h49 == _myNewVec_72_T_3[6:0] ? myVec_73 : _GEN_7282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7284 = 7'h4a == _myNewVec_72_T_3[6:0] ? myVec_74 : _GEN_7283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7285 = 7'h4b == _myNewVec_72_T_3[6:0] ? myVec_75 : _GEN_7284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7286 = 7'h4c == _myNewVec_72_T_3[6:0] ? myVec_76 : _GEN_7285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7287 = 7'h4d == _myNewVec_72_T_3[6:0] ? myVec_77 : _GEN_7286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7288 = 7'h4e == _myNewVec_72_T_3[6:0] ? myVec_78 : _GEN_7287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7289 = 7'h4f == _myNewVec_72_T_3[6:0] ? myVec_79 : _GEN_7288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7290 = 7'h50 == _myNewVec_72_T_3[6:0] ? myVec_80 : _GEN_7289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7291 = 7'h51 == _myNewVec_72_T_3[6:0] ? myVec_81 : _GEN_7290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7292 = 7'h52 == _myNewVec_72_T_3[6:0] ? myVec_82 : _GEN_7291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7293 = 7'h53 == _myNewVec_72_T_3[6:0] ? myVec_83 : _GEN_7292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7294 = 7'h54 == _myNewVec_72_T_3[6:0] ? myVec_84 : _GEN_7293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7295 = 7'h55 == _myNewVec_72_T_3[6:0] ? myVec_85 : _GEN_7294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7296 = 7'h56 == _myNewVec_72_T_3[6:0] ? myVec_86 : _GEN_7295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7297 = 7'h57 == _myNewVec_72_T_3[6:0] ? myVec_87 : _GEN_7296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7298 = 7'h58 == _myNewVec_72_T_3[6:0] ? myVec_88 : _GEN_7297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7299 = 7'h59 == _myNewVec_72_T_3[6:0] ? myVec_89 : _GEN_7298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7300 = 7'h5a == _myNewVec_72_T_3[6:0] ? myVec_90 : _GEN_7299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7301 = 7'h5b == _myNewVec_72_T_3[6:0] ? myVec_91 : _GEN_7300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7302 = 7'h5c == _myNewVec_72_T_3[6:0] ? myVec_92 : _GEN_7301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7303 = 7'h5d == _myNewVec_72_T_3[6:0] ? myVec_93 : _GEN_7302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7304 = 7'h5e == _myNewVec_72_T_3[6:0] ? myVec_94 : _GEN_7303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7305 = 7'h5f == _myNewVec_72_T_3[6:0] ? myVec_95 : _GEN_7304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7306 = 7'h60 == _myNewVec_72_T_3[6:0] ? myVec_96 : _GEN_7305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7307 = 7'h61 == _myNewVec_72_T_3[6:0] ? myVec_97 : _GEN_7306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7308 = 7'h62 == _myNewVec_72_T_3[6:0] ? myVec_98 : _GEN_7307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7309 = 7'h63 == _myNewVec_72_T_3[6:0] ? myVec_99 : _GEN_7308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7310 = 7'h64 == _myNewVec_72_T_3[6:0] ? myVec_100 : _GEN_7309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7311 = 7'h65 == _myNewVec_72_T_3[6:0] ? myVec_101 : _GEN_7310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7312 = 7'h66 == _myNewVec_72_T_3[6:0] ? myVec_102 : _GEN_7311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7313 = 7'h67 == _myNewVec_72_T_3[6:0] ? myVec_103 : _GEN_7312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7314 = 7'h68 == _myNewVec_72_T_3[6:0] ? myVec_104 : _GEN_7313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7315 = 7'h69 == _myNewVec_72_T_3[6:0] ? myVec_105 : _GEN_7314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7316 = 7'h6a == _myNewVec_72_T_3[6:0] ? myVec_106 : _GEN_7315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7317 = 7'h6b == _myNewVec_72_T_3[6:0] ? myVec_107 : _GEN_7316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7318 = 7'h6c == _myNewVec_72_T_3[6:0] ? myVec_108 : _GEN_7317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7319 = 7'h6d == _myNewVec_72_T_3[6:0] ? myVec_109 : _GEN_7318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7320 = 7'h6e == _myNewVec_72_T_3[6:0] ? myVec_110 : _GEN_7319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7321 = 7'h6f == _myNewVec_72_T_3[6:0] ? myVec_111 : _GEN_7320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7322 = 7'h70 == _myNewVec_72_T_3[6:0] ? myVec_112 : _GEN_7321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7323 = 7'h71 == _myNewVec_72_T_3[6:0] ? myVec_113 : _GEN_7322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7324 = 7'h72 == _myNewVec_72_T_3[6:0] ? myVec_114 : _GEN_7323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7325 = 7'h73 == _myNewVec_72_T_3[6:0] ? myVec_115 : _GEN_7324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7326 = 7'h74 == _myNewVec_72_T_3[6:0] ? myVec_116 : _GEN_7325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7327 = 7'h75 == _myNewVec_72_T_3[6:0] ? myVec_117 : _GEN_7326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7328 = 7'h76 == _myNewVec_72_T_3[6:0] ? myVec_118 : _GEN_7327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7329 = 7'h77 == _myNewVec_72_T_3[6:0] ? myVec_119 : _GEN_7328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7330 = 7'h78 == _myNewVec_72_T_3[6:0] ? myVec_120 : _GEN_7329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7331 = 7'h79 == _myNewVec_72_T_3[6:0] ? myVec_121 : _GEN_7330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7332 = 7'h7a == _myNewVec_72_T_3[6:0] ? myVec_122 : _GEN_7331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7333 = 7'h7b == _myNewVec_72_T_3[6:0] ? myVec_123 : _GEN_7332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7334 = 7'h7c == _myNewVec_72_T_3[6:0] ? myVec_124 : _GEN_7333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7335 = 7'h7d == _myNewVec_72_T_3[6:0] ? myVec_125 : _GEN_7334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7336 = 7'h7e == _myNewVec_72_T_3[6:0] ? myVec_126 : _GEN_7335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_72 = 7'h7f == _myNewVec_72_T_3[6:0] ? myVec_127 : _GEN_7336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_71_T_3 = _myNewVec_127_T_1 + 16'h38; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_7339 = 7'h1 == _myNewVec_71_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7340 = 7'h2 == _myNewVec_71_T_3[6:0] ? myVec_2 : _GEN_7339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7341 = 7'h3 == _myNewVec_71_T_3[6:0] ? myVec_3 : _GEN_7340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7342 = 7'h4 == _myNewVec_71_T_3[6:0] ? myVec_4 : _GEN_7341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7343 = 7'h5 == _myNewVec_71_T_3[6:0] ? myVec_5 : _GEN_7342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7344 = 7'h6 == _myNewVec_71_T_3[6:0] ? myVec_6 : _GEN_7343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7345 = 7'h7 == _myNewVec_71_T_3[6:0] ? myVec_7 : _GEN_7344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7346 = 7'h8 == _myNewVec_71_T_3[6:0] ? myVec_8 : _GEN_7345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7347 = 7'h9 == _myNewVec_71_T_3[6:0] ? myVec_9 : _GEN_7346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7348 = 7'ha == _myNewVec_71_T_3[6:0] ? myVec_10 : _GEN_7347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7349 = 7'hb == _myNewVec_71_T_3[6:0] ? myVec_11 : _GEN_7348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7350 = 7'hc == _myNewVec_71_T_3[6:0] ? myVec_12 : _GEN_7349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7351 = 7'hd == _myNewVec_71_T_3[6:0] ? myVec_13 : _GEN_7350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7352 = 7'he == _myNewVec_71_T_3[6:0] ? myVec_14 : _GEN_7351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7353 = 7'hf == _myNewVec_71_T_3[6:0] ? myVec_15 : _GEN_7352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7354 = 7'h10 == _myNewVec_71_T_3[6:0] ? myVec_16 : _GEN_7353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7355 = 7'h11 == _myNewVec_71_T_3[6:0] ? myVec_17 : _GEN_7354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7356 = 7'h12 == _myNewVec_71_T_3[6:0] ? myVec_18 : _GEN_7355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7357 = 7'h13 == _myNewVec_71_T_3[6:0] ? myVec_19 : _GEN_7356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7358 = 7'h14 == _myNewVec_71_T_3[6:0] ? myVec_20 : _GEN_7357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7359 = 7'h15 == _myNewVec_71_T_3[6:0] ? myVec_21 : _GEN_7358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7360 = 7'h16 == _myNewVec_71_T_3[6:0] ? myVec_22 : _GEN_7359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7361 = 7'h17 == _myNewVec_71_T_3[6:0] ? myVec_23 : _GEN_7360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7362 = 7'h18 == _myNewVec_71_T_3[6:0] ? myVec_24 : _GEN_7361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7363 = 7'h19 == _myNewVec_71_T_3[6:0] ? myVec_25 : _GEN_7362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7364 = 7'h1a == _myNewVec_71_T_3[6:0] ? myVec_26 : _GEN_7363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7365 = 7'h1b == _myNewVec_71_T_3[6:0] ? myVec_27 : _GEN_7364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7366 = 7'h1c == _myNewVec_71_T_3[6:0] ? myVec_28 : _GEN_7365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7367 = 7'h1d == _myNewVec_71_T_3[6:0] ? myVec_29 : _GEN_7366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7368 = 7'h1e == _myNewVec_71_T_3[6:0] ? myVec_30 : _GEN_7367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7369 = 7'h1f == _myNewVec_71_T_3[6:0] ? myVec_31 : _GEN_7368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7370 = 7'h20 == _myNewVec_71_T_3[6:0] ? myVec_32 : _GEN_7369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7371 = 7'h21 == _myNewVec_71_T_3[6:0] ? myVec_33 : _GEN_7370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7372 = 7'h22 == _myNewVec_71_T_3[6:0] ? myVec_34 : _GEN_7371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7373 = 7'h23 == _myNewVec_71_T_3[6:0] ? myVec_35 : _GEN_7372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7374 = 7'h24 == _myNewVec_71_T_3[6:0] ? myVec_36 : _GEN_7373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7375 = 7'h25 == _myNewVec_71_T_3[6:0] ? myVec_37 : _GEN_7374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7376 = 7'h26 == _myNewVec_71_T_3[6:0] ? myVec_38 : _GEN_7375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7377 = 7'h27 == _myNewVec_71_T_3[6:0] ? myVec_39 : _GEN_7376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7378 = 7'h28 == _myNewVec_71_T_3[6:0] ? myVec_40 : _GEN_7377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7379 = 7'h29 == _myNewVec_71_T_3[6:0] ? myVec_41 : _GEN_7378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7380 = 7'h2a == _myNewVec_71_T_3[6:0] ? myVec_42 : _GEN_7379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7381 = 7'h2b == _myNewVec_71_T_3[6:0] ? myVec_43 : _GEN_7380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7382 = 7'h2c == _myNewVec_71_T_3[6:0] ? myVec_44 : _GEN_7381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7383 = 7'h2d == _myNewVec_71_T_3[6:0] ? myVec_45 : _GEN_7382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7384 = 7'h2e == _myNewVec_71_T_3[6:0] ? myVec_46 : _GEN_7383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7385 = 7'h2f == _myNewVec_71_T_3[6:0] ? myVec_47 : _GEN_7384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7386 = 7'h30 == _myNewVec_71_T_3[6:0] ? myVec_48 : _GEN_7385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7387 = 7'h31 == _myNewVec_71_T_3[6:0] ? myVec_49 : _GEN_7386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7388 = 7'h32 == _myNewVec_71_T_3[6:0] ? myVec_50 : _GEN_7387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7389 = 7'h33 == _myNewVec_71_T_3[6:0] ? myVec_51 : _GEN_7388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7390 = 7'h34 == _myNewVec_71_T_3[6:0] ? myVec_52 : _GEN_7389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7391 = 7'h35 == _myNewVec_71_T_3[6:0] ? myVec_53 : _GEN_7390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7392 = 7'h36 == _myNewVec_71_T_3[6:0] ? myVec_54 : _GEN_7391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7393 = 7'h37 == _myNewVec_71_T_3[6:0] ? myVec_55 : _GEN_7392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7394 = 7'h38 == _myNewVec_71_T_3[6:0] ? myVec_56 : _GEN_7393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7395 = 7'h39 == _myNewVec_71_T_3[6:0] ? myVec_57 : _GEN_7394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7396 = 7'h3a == _myNewVec_71_T_3[6:0] ? myVec_58 : _GEN_7395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7397 = 7'h3b == _myNewVec_71_T_3[6:0] ? myVec_59 : _GEN_7396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7398 = 7'h3c == _myNewVec_71_T_3[6:0] ? myVec_60 : _GEN_7397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7399 = 7'h3d == _myNewVec_71_T_3[6:0] ? myVec_61 : _GEN_7398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7400 = 7'h3e == _myNewVec_71_T_3[6:0] ? myVec_62 : _GEN_7399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7401 = 7'h3f == _myNewVec_71_T_3[6:0] ? myVec_63 : _GEN_7400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7402 = 7'h40 == _myNewVec_71_T_3[6:0] ? myVec_64 : _GEN_7401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7403 = 7'h41 == _myNewVec_71_T_3[6:0] ? myVec_65 : _GEN_7402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7404 = 7'h42 == _myNewVec_71_T_3[6:0] ? myVec_66 : _GEN_7403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7405 = 7'h43 == _myNewVec_71_T_3[6:0] ? myVec_67 : _GEN_7404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7406 = 7'h44 == _myNewVec_71_T_3[6:0] ? myVec_68 : _GEN_7405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7407 = 7'h45 == _myNewVec_71_T_3[6:0] ? myVec_69 : _GEN_7406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7408 = 7'h46 == _myNewVec_71_T_3[6:0] ? myVec_70 : _GEN_7407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7409 = 7'h47 == _myNewVec_71_T_3[6:0] ? myVec_71 : _GEN_7408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7410 = 7'h48 == _myNewVec_71_T_3[6:0] ? myVec_72 : _GEN_7409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7411 = 7'h49 == _myNewVec_71_T_3[6:0] ? myVec_73 : _GEN_7410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7412 = 7'h4a == _myNewVec_71_T_3[6:0] ? myVec_74 : _GEN_7411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7413 = 7'h4b == _myNewVec_71_T_3[6:0] ? myVec_75 : _GEN_7412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7414 = 7'h4c == _myNewVec_71_T_3[6:0] ? myVec_76 : _GEN_7413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7415 = 7'h4d == _myNewVec_71_T_3[6:0] ? myVec_77 : _GEN_7414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7416 = 7'h4e == _myNewVec_71_T_3[6:0] ? myVec_78 : _GEN_7415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7417 = 7'h4f == _myNewVec_71_T_3[6:0] ? myVec_79 : _GEN_7416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7418 = 7'h50 == _myNewVec_71_T_3[6:0] ? myVec_80 : _GEN_7417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7419 = 7'h51 == _myNewVec_71_T_3[6:0] ? myVec_81 : _GEN_7418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7420 = 7'h52 == _myNewVec_71_T_3[6:0] ? myVec_82 : _GEN_7419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7421 = 7'h53 == _myNewVec_71_T_3[6:0] ? myVec_83 : _GEN_7420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7422 = 7'h54 == _myNewVec_71_T_3[6:0] ? myVec_84 : _GEN_7421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7423 = 7'h55 == _myNewVec_71_T_3[6:0] ? myVec_85 : _GEN_7422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7424 = 7'h56 == _myNewVec_71_T_3[6:0] ? myVec_86 : _GEN_7423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7425 = 7'h57 == _myNewVec_71_T_3[6:0] ? myVec_87 : _GEN_7424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7426 = 7'h58 == _myNewVec_71_T_3[6:0] ? myVec_88 : _GEN_7425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7427 = 7'h59 == _myNewVec_71_T_3[6:0] ? myVec_89 : _GEN_7426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7428 = 7'h5a == _myNewVec_71_T_3[6:0] ? myVec_90 : _GEN_7427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7429 = 7'h5b == _myNewVec_71_T_3[6:0] ? myVec_91 : _GEN_7428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7430 = 7'h5c == _myNewVec_71_T_3[6:0] ? myVec_92 : _GEN_7429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7431 = 7'h5d == _myNewVec_71_T_3[6:0] ? myVec_93 : _GEN_7430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7432 = 7'h5e == _myNewVec_71_T_3[6:0] ? myVec_94 : _GEN_7431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7433 = 7'h5f == _myNewVec_71_T_3[6:0] ? myVec_95 : _GEN_7432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7434 = 7'h60 == _myNewVec_71_T_3[6:0] ? myVec_96 : _GEN_7433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7435 = 7'h61 == _myNewVec_71_T_3[6:0] ? myVec_97 : _GEN_7434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7436 = 7'h62 == _myNewVec_71_T_3[6:0] ? myVec_98 : _GEN_7435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7437 = 7'h63 == _myNewVec_71_T_3[6:0] ? myVec_99 : _GEN_7436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7438 = 7'h64 == _myNewVec_71_T_3[6:0] ? myVec_100 : _GEN_7437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7439 = 7'h65 == _myNewVec_71_T_3[6:0] ? myVec_101 : _GEN_7438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7440 = 7'h66 == _myNewVec_71_T_3[6:0] ? myVec_102 : _GEN_7439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7441 = 7'h67 == _myNewVec_71_T_3[6:0] ? myVec_103 : _GEN_7440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7442 = 7'h68 == _myNewVec_71_T_3[6:0] ? myVec_104 : _GEN_7441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7443 = 7'h69 == _myNewVec_71_T_3[6:0] ? myVec_105 : _GEN_7442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7444 = 7'h6a == _myNewVec_71_T_3[6:0] ? myVec_106 : _GEN_7443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7445 = 7'h6b == _myNewVec_71_T_3[6:0] ? myVec_107 : _GEN_7444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7446 = 7'h6c == _myNewVec_71_T_3[6:0] ? myVec_108 : _GEN_7445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7447 = 7'h6d == _myNewVec_71_T_3[6:0] ? myVec_109 : _GEN_7446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7448 = 7'h6e == _myNewVec_71_T_3[6:0] ? myVec_110 : _GEN_7447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7449 = 7'h6f == _myNewVec_71_T_3[6:0] ? myVec_111 : _GEN_7448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7450 = 7'h70 == _myNewVec_71_T_3[6:0] ? myVec_112 : _GEN_7449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7451 = 7'h71 == _myNewVec_71_T_3[6:0] ? myVec_113 : _GEN_7450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7452 = 7'h72 == _myNewVec_71_T_3[6:0] ? myVec_114 : _GEN_7451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7453 = 7'h73 == _myNewVec_71_T_3[6:0] ? myVec_115 : _GEN_7452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7454 = 7'h74 == _myNewVec_71_T_3[6:0] ? myVec_116 : _GEN_7453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7455 = 7'h75 == _myNewVec_71_T_3[6:0] ? myVec_117 : _GEN_7454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7456 = 7'h76 == _myNewVec_71_T_3[6:0] ? myVec_118 : _GEN_7455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7457 = 7'h77 == _myNewVec_71_T_3[6:0] ? myVec_119 : _GEN_7456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7458 = 7'h78 == _myNewVec_71_T_3[6:0] ? myVec_120 : _GEN_7457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7459 = 7'h79 == _myNewVec_71_T_3[6:0] ? myVec_121 : _GEN_7458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7460 = 7'h7a == _myNewVec_71_T_3[6:0] ? myVec_122 : _GEN_7459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7461 = 7'h7b == _myNewVec_71_T_3[6:0] ? myVec_123 : _GEN_7460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7462 = 7'h7c == _myNewVec_71_T_3[6:0] ? myVec_124 : _GEN_7461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7463 = 7'h7d == _myNewVec_71_T_3[6:0] ? myVec_125 : _GEN_7462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7464 = 7'h7e == _myNewVec_71_T_3[6:0] ? myVec_126 : _GEN_7463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_71 = 7'h7f == _myNewVec_71_T_3[6:0] ? myVec_127 : _GEN_7464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_70_T_3 = _myNewVec_127_T_1 + 16'h39; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_7467 = 7'h1 == _myNewVec_70_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7468 = 7'h2 == _myNewVec_70_T_3[6:0] ? myVec_2 : _GEN_7467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7469 = 7'h3 == _myNewVec_70_T_3[6:0] ? myVec_3 : _GEN_7468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7470 = 7'h4 == _myNewVec_70_T_3[6:0] ? myVec_4 : _GEN_7469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7471 = 7'h5 == _myNewVec_70_T_3[6:0] ? myVec_5 : _GEN_7470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7472 = 7'h6 == _myNewVec_70_T_3[6:0] ? myVec_6 : _GEN_7471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7473 = 7'h7 == _myNewVec_70_T_3[6:0] ? myVec_7 : _GEN_7472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7474 = 7'h8 == _myNewVec_70_T_3[6:0] ? myVec_8 : _GEN_7473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7475 = 7'h9 == _myNewVec_70_T_3[6:0] ? myVec_9 : _GEN_7474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7476 = 7'ha == _myNewVec_70_T_3[6:0] ? myVec_10 : _GEN_7475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7477 = 7'hb == _myNewVec_70_T_3[6:0] ? myVec_11 : _GEN_7476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7478 = 7'hc == _myNewVec_70_T_3[6:0] ? myVec_12 : _GEN_7477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7479 = 7'hd == _myNewVec_70_T_3[6:0] ? myVec_13 : _GEN_7478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7480 = 7'he == _myNewVec_70_T_3[6:0] ? myVec_14 : _GEN_7479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7481 = 7'hf == _myNewVec_70_T_3[6:0] ? myVec_15 : _GEN_7480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7482 = 7'h10 == _myNewVec_70_T_3[6:0] ? myVec_16 : _GEN_7481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7483 = 7'h11 == _myNewVec_70_T_3[6:0] ? myVec_17 : _GEN_7482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7484 = 7'h12 == _myNewVec_70_T_3[6:0] ? myVec_18 : _GEN_7483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7485 = 7'h13 == _myNewVec_70_T_3[6:0] ? myVec_19 : _GEN_7484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7486 = 7'h14 == _myNewVec_70_T_3[6:0] ? myVec_20 : _GEN_7485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7487 = 7'h15 == _myNewVec_70_T_3[6:0] ? myVec_21 : _GEN_7486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7488 = 7'h16 == _myNewVec_70_T_3[6:0] ? myVec_22 : _GEN_7487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7489 = 7'h17 == _myNewVec_70_T_3[6:0] ? myVec_23 : _GEN_7488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7490 = 7'h18 == _myNewVec_70_T_3[6:0] ? myVec_24 : _GEN_7489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7491 = 7'h19 == _myNewVec_70_T_3[6:0] ? myVec_25 : _GEN_7490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7492 = 7'h1a == _myNewVec_70_T_3[6:0] ? myVec_26 : _GEN_7491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7493 = 7'h1b == _myNewVec_70_T_3[6:0] ? myVec_27 : _GEN_7492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7494 = 7'h1c == _myNewVec_70_T_3[6:0] ? myVec_28 : _GEN_7493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7495 = 7'h1d == _myNewVec_70_T_3[6:0] ? myVec_29 : _GEN_7494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7496 = 7'h1e == _myNewVec_70_T_3[6:0] ? myVec_30 : _GEN_7495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7497 = 7'h1f == _myNewVec_70_T_3[6:0] ? myVec_31 : _GEN_7496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7498 = 7'h20 == _myNewVec_70_T_3[6:0] ? myVec_32 : _GEN_7497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7499 = 7'h21 == _myNewVec_70_T_3[6:0] ? myVec_33 : _GEN_7498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7500 = 7'h22 == _myNewVec_70_T_3[6:0] ? myVec_34 : _GEN_7499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7501 = 7'h23 == _myNewVec_70_T_3[6:0] ? myVec_35 : _GEN_7500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7502 = 7'h24 == _myNewVec_70_T_3[6:0] ? myVec_36 : _GEN_7501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7503 = 7'h25 == _myNewVec_70_T_3[6:0] ? myVec_37 : _GEN_7502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7504 = 7'h26 == _myNewVec_70_T_3[6:0] ? myVec_38 : _GEN_7503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7505 = 7'h27 == _myNewVec_70_T_3[6:0] ? myVec_39 : _GEN_7504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7506 = 7'h28 == _myNewVec_70_T_3[6:0] ? myVec_40 : _GEN_7505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7507 = 7'h29 == _myNewVec_70_T_3[6:0] ? myVec_41 : _GEN_7506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7508 = 7'h2a == _myNewVec_70_T_3[6:0] ? myVec_42 : _GEN_7507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7509 = 7'h2b == _myNewVec_70_T_3[6:0] ? myVec_43 : _GEN_7508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7510 = 7'h2c == _myNewVec_70_T_3[6:0] ? myVec_44 : _GEN_7509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7511 = 7'h2d == _myNewVec_70_T_3[6:0] ? myVec_45 : _GEN_7510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7512 = 7'h2e == _myNewVec_70_T_3[6:0] ? myVec_46 : _GEN_7511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7513 = 7'h2f == _myNewVec_70_T_3[6:0] ? myVec_47 : _GEN_7512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7514 = 7'h30 == _myNewVec_70_T_3[6:0] ? myVec_48 : _GEN_7513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7515 = 7'h31 == _myNewVec_70_T_3[6:0] ? myVec_49 : _GEN_7514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7516 = 7'h32 == _myNewVec_70_T_3[6:0] ? myVec_50 : _GEN_7515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7517 = 7'h33 == _myNewVec_70_T_3[6:0] ? myVec_51 : _GEN_7516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7518 = 7'h34 == _myNewVec_70_T_3[6:0] ? myVec_52 : _GEN_7517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7519 = 7'h35 == _myNewVec_70_T_3[6:0] ? myVec_53 : _GEN_7518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7520 = 7'h36 == _myNewVec_70_T_3[6:0] ? myVec_54 : _GEN_7519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7521 = 7'h37 == _myNewVec_70_T_3[6:0] ? myVec_55 : _GEN_7520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7522 = 7'h38 == _myNewVec_70_T_3[6:0] ? myVec_56 : _GEN_7521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7523 = 7'h39 == _myNewVec_70_T_3[6:0] ? myVec_57 : _GEN_7522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7524 = 7'h3a == _myNewVec_70_T_3[6:0] ? myVec_58 : _GEN_7523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7525 = 7'h3b == _myNewVec_70_T_3[6:0] ? myVec_59 : _GEN_7524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7526 = 7'h3c == _myNewVec_70_T_3[6:0] ? myVec_60 : _GEN_7525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7527 = 7'h3d == _myNewVec_70_T_3[6:0] ? myVec_61 : _GEN_7526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7528 = 7'h3e == _myNewVec_70_T_3[6:0] ? myVec_62 : _GEN_7527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7529 = 7'h3f == _myNewVec_70_T_3[6:0] ? myVec_63 : _GEN_7528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7530 = 7'h40 == _myNewVec_70_T_3[6:0] ? myVec_64 : _GEN_7529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7531 = 7'h41 == _myNewVec_70_T_3[6:0] ? myVec_65 : _GEN_7530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7532 = 7'h42 == _myNewVec_70_T_3[6:0] ? myVec_66 : _GEN_7531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7533 = 7'h43 == _myNewVec_70_T_3[6:0] ? myVec_67 : _GEN_7532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7534 = 7'h44 == _myNewVec_70_T_3[6:0] ? myVec_68 : _GEN_7533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7535 = 7'h45 == _myNewVec_70_T_3[6:0] ? myVec_69 : _GEN_7534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7536 = 7'h46 == _myNewVec_70_T_3[6:0] ? myVec_70 : _GEN_7535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7537 = 7'h47 == _myNewVec_70_T_3[6:0] ? myVec_71 : _GEN_7536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7538 = 7'h48 == _myNewVec_70_T_3[6:0] ? myVec_72 : _GEN_7537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7539 = 7'h49 == _myNewVec_70_T_3[6:0] ? myVec_73 : _GEN_7538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7540 = 7'h4a == _myNewVec_70_T_3[6:0] ? myVec_74 : _GEN_7539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7541 = 7'h4b == _myNewVec_70_T_3[6:0] ? myVec_75 : _GEN_7540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7542 = 7'h4c == _myNewVec_70_T_3[6:0] ? myVec_76 : _GEN_7541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7543 = 7'h4d == _myNewVec_70_T_3[6:0] ? myVec_77 : _GEN_7542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7544 = 7'h4e == _myNewVec_70_T_3[6:0] ? myVec_78 : _GEN_7543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7545 = 7'h4f == _myNewVec_70_T_3[6:0] ? myVec_79 : _GEN_7544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7546 = 7'h50 == _myNewVec_70_T_3[6:0] ? myVec_80 : _GEN_7545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7547 = 7'h51 == _myNewVec_70_T_3[6:0] ? myVec_81 : _GEN_7546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7548 = 7'h52 == _myNewVec_70_T_3[6:0] ? myVec_82 : _GEN_7547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7549 = 7'h53 == _myNewVec_70_T_3[6:0] ? myVec_83 : _GEN_7548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7550 = 7'h54 == _myNewVec_70_T_3[6:0] ? myVec_84 : _GEN_7549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7551 = 7'h55 == _myNewVec_70_T_3[6:0] ? myVec_85 : _GEN_7550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7552 = 7'h56 == _myNewVec_70_T_3[6:0] ? myVec_86 : _GEN_7551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7553 = 7'h57 == _myNewVec_70_T_3[6:0] ? myVec_87 : _GEN_7552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7554 = 7'h58 == _myNewVec_70_T_3[6:0] ? myVec_88 : _GEN_7553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7555 = 7'h59 == _myNewVec_70_T_3[6:0] ? myVec_89 : _GEN_7554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7556 = 7'h5a == _myNewVec_70_T_3[6:0] ? myVec_90 : _GEN_7555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7557 = 7'h5b == _myNewVec_70_T_3[6:0] ? myVec_91 : _GEN_7556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7558 = 7'h5c == _myNewVec_70_T_3[6:0] ? myVec_92 : _GEN_7557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7559 = 7'h5d == _myNewVec_70_T_3[6:0] ? myVec_93 : _GEN_7558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7560 = 7'h5e == _myNewVec_70_T_3[6:0] ? myVec_94 : _GEN_7559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7561 = 7'h5f == _myNewVec_70_T_3[6:0] ? myVec_95 : _GEN_7560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7562 = 7'h60 == _myNewVec_70_T_3[6:0] ? myVec_96 : _GEN_7561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7563 = 7'h61 == _myNewVec_70_T_3[6:0] ? myVec_97 : _GEN_7562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7564 = 7'h62 == _myNewVec_70_T_3[6:0] ? myVec_98 : _GEN_7563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7565 = 7'h63 == _myNewVec_70_T_3[6:0] ? myVec_99 : _GEN_7564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7566 = 7'h64 == _myNewVec_70_T_3[6:0] ? myVec_100 : _GEN_7565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7567 = 7'h65 == _myNewVec_70_T_3[6:0] ? myVec_101 : _GEN_7566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7568 = 7'h66 == _myNewVec_70_T_3[6:0] ? myVec_102 : _GEN_7567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7569 = 7'h67 == _myNewVec_70_T_3[6:0] ? myVec_103 : _GEN_7568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7570 = 7'h68 == _myNewVec_70_T_3[6:0] ? myVec_104 : _GEN_7569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7571 = 7'h69 == _myNewVec_70_T_3[6:0] ? myVec_105 : _GEN_7570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7572 = 7'h6a == _myNewVec_70_T_3[6:0] ? myVec_106 : _GEN_7571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7573 = 7'h6b == _myNewVec_70_T_3[6:0] ? myVec_107 : _GEN_7572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7574 = 7'h6c == _myNewVec_70_T_3[6:0] ? myVec_108 : _GEN_7573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7575 = 7'h6d == _myNewVec_70_T_3[6:0] ? myVec_109 : _GEN_7574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7576 = 7'h6e == _myNewVec_70_T_3[6:0] ? myVec_110 : _GEN_7575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7577 = 7'h6f == _myNewVec_70_T_3[6:0] ? myVec_111 : _GEN_7576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7578 = 7'h70 == _myNewVec_70_T_3[6:0] ? myVec_112 : _GEN_7577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7579 = 7'h71 == _myNewVec_70_T_3[6:0] ? myVec_113 : _GEN_7578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7580 = 7'h72 == _myNewVec_70_T_3[6:0] ? myVec_114 : _GEN_7579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7581 = 7'h73 == _myNewVec_70_T_3[6:0] ? myVec_115 : _GEN_7580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7582 = 7'h74 == _myNewVec_70_T_3[6:0] ? myVec_116 : _GEN_7581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7583 = 7'h75 == _myNewVec_70_T_3[6:0] ? myVec_117 : _GEN_7582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7584 = 7'h76 == _myNewVec_70_T_3[6:0] ? myVec_118 : _GEN_7583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7585 = 7'h77 == _myNewVec_70_T_3[6:0] ? myVec_119 : _GEN_7584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7586 = 7'h78 == _myNewVec_70_T_3[6:0] ? myVec_120 : _GEN_7585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7587 = 7'h79 == _myNewVec_70_T_3[6:0] ? myVec_121 : _GEN_7586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7588 = 7'h7a == _myNewVec_70_T_3[6:0] ? myVec_122 : _GEN_7587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7589 = 7'h7b == _myNewVec_70_T_3[6:0] ? myVec_123 : _GEN_7588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7590 = 7'h7c == _myNewVec_70_T_3[6:0] ? myVec_124 : _GEN_7589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7591 = 7'h7d == _myNewVec_70_T_3[6:0] ? myVec_125 : _GEN_7590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7592 = 7'h7e == _myNewVec_70_T_3[6:0] ? myVec_126 : _GEN_7591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_70 = 7'h7f == _myNewVec_70_T_3[6:0] ? myVec_127 : _GEN_7592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_69_T_3 = _myNewVec_127_T_1 + 16'h3a; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_7595 = 7'h1 == _myNewVec_69_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7596 = 7'h2 == _myNewVec_69_T_3[6:0] ? myVec_2 : _GEN_7595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7597 = 7'h3 == _myNewVec_69_T_3[6:0] ? myVec_3 : _GEN_7596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7598 = 7'h4 == _myNewVec_69_T_3[6:0] ? myVec_4 : _GEN_7597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7599 = 7'h5 == _myNewVec_69_T_3[6:0] ? myVec_5 : _GEN_7598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7600 = 7'h6 == _myNewVec_69_T_3[6:0] ? myVec_6 : _GEN_7599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7601 = 7'h7 == _myNewVec_69_T_3[6:0] ? myVec_7 : _GEN_7600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7602 = 7'h8 == _myNewVec_69_T_3[6:0] ? myVec_8 : _GEN_7601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7603 = 7'h9 == _myNewVec_69_T_3[6:0] ? myVec_9 : _GEN_7602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7604 = 7'ha == _myNewVec_69_T_3[6:0] ? myVec_10 : _GEN_7603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7605 = 7'hb == _myNewVec_69_T_3[6:0] ? myVec_11 : _GEN_7604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7606 = 7'hc == _myNewVec_69_T_3[6:0] ? myVec_12 : _GEN_7605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7607 = 7'hd == _myNewVec_69_T_3[6:0] ? myVec_13 : _GEN_7606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7608 = 7'he == _myNewVec_69_T_3[6:0] ? myVec_14 : _GEN_7607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7609 = 7'hf == _myNewVec_69_T_3[6:0] ? myVec_15 : _GEN_7608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7610 = 7'h10 == _myNewVec_69_T_3[6:0] ? myVec_16 : _GEN_7609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7611 = 7'h11 == _myNewVec_69_T_3[6:0] ? myVec_17 : _GEN_7610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7612 = 7'h12 == _myNewVec_69_T_3[6:0] ? myVec_18 : _GEN_7611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7613 = 7'h13 == _myNewVec_69_T_3[6:0] ? myVec_19 : _GEN_7612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7614 = 7'h14 == _myNewVec_69_T_3[6:0] ? myVec_20 : _GEN_7613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7615 = 7'h15 == _myNewVec_69_T_3[6:0] ? myVec_21 : _GEN_7614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7616 = 7'h16 == _myNewVec_69_T_3[6:0] ? myVec_22 : _GEN_7615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7617 = 7'h17 == _myNewVec_69_T_3[6:0] ? myVec_23 : _GEN_7616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7618 = 7'h18 == _myNewVec_69_T_3[6:0] ? myVec_24 : _GEN_7617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7619 = 7'h19 == _myNewVec_69_T_3[6:0] ? myVec_25 : _GEN_7618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7620 = 7'h1a == _myNewVec_69_T_3[6:0] ? myVec_26 : _GEN_7619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7621 = 7'h1b == _myNewVec_69_T_3[6:0] ? myVec_27 : _GEN_7620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7622 = 7'h1c == _myNewVec_69_T_3[6:0] ? myVec_28 : _GEN_7621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7623 = 7'h1d == _myNewVec_69_T_3[6:0] ? myVec_29 : _GEN_7622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7624 = 7'h1e == _myNewVec_69_T_3[6:0] ? myVec_30 : _GEN_7623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7625 = 7'h1f == _myNewVec_69_T_3[6:0] ? myVec_31 : _GEN_7624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7626 = 7'h20 == _myNewVec_69_T_3[6:0] ? myVec_32 : _GEN_7625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7627 = 7'h21 == _myNewVec_69_T_3[6:0] ? myVec_33 : _GEN_7626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7628 = 7'h22 == _myNewVec_69_T_3[6:0] ? myVec_34 : _GEN_7627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7629 = 7'h23 == _myNewVec_69_T_3[6:0] ? myVec_35 : _GEN_7628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7630 = 7'h24 == _myNewVec_69_T_3[6:0] ? myVec_36 : _GEN_7629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7631 = 7'h25 == _myNewVec_69_T_3[6:0] ? myVec_37 : _GEN_7630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7632 = 7'h26 == _myNewVec_69_T_3[6:0] ? myVec_38 : _GEN_7631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7633 = 7'h27 == _myNewVec_69_T_3[6:0] ? myVec_39 : _GEN_7632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7634 = 7'h28 == _myNewVec_69_T_3[6:0] ? myVec_40 : _GEN_7633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7635 = 7'h29 == _myNewVec_69_T_3[6:0] ? myVec_41 : _GEN_7634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7636 = 7'h2a == _myNewVec_69_T_3[6:0] ? myVec_42 : _GEN_7635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7637 = 7'h2b == _myNewVec_69_T_3[6:0] ? myVec_43 : _GEN_7636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7638 = 7'h2c == _myNewVec_69_T_3[6:0] ? myVec_44 : _GEN_7637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7639 = 7'h2d == _myNewVec_69_T_3[6:0] ? myVec_45 : _GEN_7638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7640 = 7'h2e == _myNewVec_69_T_3[6:0] ? myVec_46 : _GEN_7639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7641 = 7'h2f == _myNewVec_69_T_3[6:0] ? myVec_47 : _GEN_7640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7642 = 7'h30 == _myNewVec_69_T_3[6:0] ? myVec_48 : _GEN_7641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7643 = 7'h31 == _myNewVec_69_T_3[6:0] ? myVec_49 : _GEN_7642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7644 = 7'h32 == _myNewVec_69_T_3[6:0] ? myVec_50 : _GEN_7643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7645 = 7'h33 == _myNewVec_69_T_3[6:0] ? myVec_51 : _GEN_7644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7646 = 7'h34 == _myNewVec_69_T_3[6:0] ? myVec_52 : _GEN_7645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7647 = 7'h35 == _myNewVec_69_T_3[6:0] ? myVec_53 : _GEN_7646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7648 = 7'h36 == _myNewVec_69_T_3[6:0] ? myVec_54 : _GEN_7647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7649 = 7'h37 == _myNewVec_69_T_3[6:0] ? myVec_55 : _GEN_7648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7650 = 7'h38 == _myNewVec_69_T_3[6:0] ? myVec_56 : _GEN_7649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7651 = 7'h39 == _myNewVec_69_T_3[6:0] ? myVec_57 : _GEN_7650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7652 = 7'h3a == _myNewVec_69_T_3[6:0] ? myVec_58 : _GEN_7651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7653 = 7'h3b == _myNewVec_69_T_3[6:0] ? myVec_59 : _GEN_7652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7654 = 7'h3c == _myNewVec_69_T_3[6:0] ? myVec_60 : _GEN_7653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7655 = 7'h3d == _myNewVec_69_T_3[6:0] ? myVec_61 : _GEN_7654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7656 = 7'h3e == _myNewVec_69_T_3[6:0] ? myVec_62 : _GEN_7655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7657 = 7'h3f == _myNewVec_69_T_3[6:0] ? myVec_63 : _GEN_7656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7658 = 7'h40 == _myNewVec_69_T_3[6:0] ? myVec_64 : _GEN_7657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7659 = 7'h41 == _myNewVec_69_T_3[6:0] ? myVec_65 : _GEN_7658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7660 = 7'h42 == _myNewVec_69_T_3[6:0] ? myVec_66 : _GEN_7659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7661 = 7'h43 == _myNewVec_69_T_3[6:0] ? myVec_67 : _GEN_7660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7662 = 7'h44 == _myNewVec_69_T_3[6:0] ? myVec_68 : _GEN_7661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7663 = 7'h45 == _myNewVec_69_T_3[6:0] ? myVec_69 : _GEN_7662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7664 = 7'h46 == _myNewVec_69_T_3[6:0] ? myVec_70 : _GEN_7663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7665 = 7'h47 == _myNewVec_69_T_3[6:0] ? myVec_71 : _GEN_7664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7666 = 7'h48 == _myNewVec_69_T_3[6:0] ? myVec_72 : _GEN_7665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7667 = 7'h49 == _myNewVec_69_T_3[6:0] ? myVec_73 : _GEN_7666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7668 = 7'h4a == _myNewVec_69_T_3[6:0] ? myVec_74 : _GEN_7667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7669 = 7'h4b == _myNewVec_69_T_3[6:0] ? myVec_75 : _GEN_7668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7670 = 7'h4c == _myNewVec_69_T_3[6:0] ? myVec_76 : _GEN_7669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7671 = 7'h4d == _myNewVec_69_T_3[6:0] ? myVec_77 : _GEN_7670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7672 = 7'h4e == _myNewVec_69_T_3[6:0] ? myVec_78 : _GEN_7671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7673 = 7'h4f == _myNewVec_69_T_3[6:0] ? myVec_79 : _GEN_7672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7674 = 7'h50 == _myNewVec_69_T_3[6:0] ? myVec_80 : _GEN_7673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7675 = 7'h51 == _myNewVec_69_T_3[6:0] ? myVec_81 : _GEN_7674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7676 = 7'h52 == _myNewVec_69_T_3[6:0] ? myVec_82 : _GEN_7675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7677 = 7'h53 == _myNewVec_69_T_3[6:0] ? myVec_83 : _GEN_7676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7678 = 7'h54 == _myNewVec_69_T_3[6:0] ? myVec_84 : _GEN_7677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7679 = 7'h55 == _myNewVec_69_T_3[6:0] ? myVec_85 : _GEN_7678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7680 = 7'h56 == _myNewVec_69_T_3[6:0] ? myVec_86 : _GEN_7679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7681 = 7'h57 == _myNewVec_69_T_3[6:0] ? myVec_87 : _GEN_7680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7682 = 7'h58 == _myNewVec_69_T_3[6:0] ? myVec_88 : _GEN_7681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7683 = 7'h59 == _myNewVec_69_T_3[6:0] ? myVec_89 : _GEN_7682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7684 = 7'h5a == _myNewVec_69_T_3[6:0] ? myVec_90 : _GEN_7683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7685 = 7'h5b == _myNewVec_69_T_3[6:0] ? myVec_91 : _GEN_7684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7686 = 7'h5c == _myNewVec_69_T_3[6:0] ? myVec_92 : _GEN_7685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7687 = 7'h5d == _myNewVec_69_T_3[6:0] ? myVec_93 : _GEN_7686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7688 = 7'h5e == _myNewVec_69_T_3[6:0] ? myVec_94 : _GEN_7687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7689 = 7'h5f == _myNewVec_69_T_3[6:0] ? myVec_95 : _GEN_7688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7690 = 7'h60 == _myNewVec_69_T_3[6:0] ? myVec_96 : _GEN_7689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7691 = 7'h61 == _myNewVec_69_T_3[6:0] ? myVec_97 : _GEN_7690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7692 = 7'h62 == _myNewVec_69_T_3[6:0] ? myVec_98 : _GEN_7691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7693 = 7'h63 == _myNewVec_69_T_3[6:0] ? myVec_99 : _GEN_7692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7694 = 7'h64 == _myNewVec_69_T_3[6:0] ? myVec_100 : _GEN_7693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7695 = 7'h65 == _myNewVec_69_T_3[6:0] ? myVec_101 : _GEN_7694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7696 = 7'h66 == _myNewVec_69_T_3[6:0] ? myVec_102 : _GEN_7695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7697 = 7'h67 == _myNewVec_69_T_3[6:0] ? myVec_103 : _GEN_7696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7698 = 7'h68 == _myNewVec_69_T_3[6:0] ? myVec_104 : _GEN_7697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7699 = 7'h69 == _myNewVec_69_T_3[6:0] ? myVec_105 : _GEN_7698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7700 = 7'h6a == _myNewVec_69_T_3[6:0] ? myVec_106 : _GEN_7699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7701 = 7'h6b == _myNewVec_69_T_3[6:0] ? myVec_107 : _GEN_7700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7702 = 7'h6c == _myNewVec_69_T_3[6:0] ? myVec_108 : _GEN_7701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7703 = 7'h6d == _myNewVec_69_T_3[6:0] ? myVec_109 : _GEN_7702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7704 = 7'h6e == _myNewVec_69_T_3[6:0] ? myVec_110 : _GEN_7703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7705 = 7'h6f == _myNewVec_69_T_3[6:0] ? myVec_111 : _GEN_7704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7706 = 7'h70 == _myNewVec_69_T_3[6:0] ? myVec_112 : _GEN_7705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7707 = 7'h71 == _myNewVec_69_T_3[6:0] ? myVec_113 : _GEN_7706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7708 = 7'h72 == _myNewVec_69_T_3[6:0] ? myVec_114 : _GEN_7707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7709 = 7'h73 == _myNewVec_69_T_3[6:0] ? myVec_115 : _GEN_7708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7710 = 7'h74 == _myNewVec_69_T_3[6:0] ? myVec_116 : _GEN_7709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7711 = 7'h75 == _myNewVec_69_T_3[6:0] ? myVec_117 : _GEN_7710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7712 = 7'h76 == _myNewVec_69_T_3[6:0] ? myVec_118 : _GEN_7711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7713 = 7'h77 == _myNewVec_69_T_3[6:0] ? myVec_119 : _GEN_7712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7714 = 7'h78 == _myNewVec_69_T_3[6:0] ? myVec_120 : _GEN_7713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7715 = 7'h79 == _myNewVec_69_T_3[6:0] ? myVec_121 : _GEN_7714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7716 = 7'h7a == _myNewVec_69_T_3[6:0] ? myVec_122 : _GEN_7715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7717 = 7'h7b == _myNewVec_69_T_3[6:0] ? myVec_123 : _GEN_7716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7718 = 7'h7c == _myNewVec_69_T_3[6:0] ? myVec_124 : _GEN_7717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7719 = 7'h7d == _myNewVec_69_T_3[6:0] ? myVec_125 : _GEN_7718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7720 = 7'h7e == _myNewVec_69_T_3[6:0] ? myVec_126 : _GEN_7719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_69 = 7'h7f == _myNewVec_69_T_3[6:0] ? myVec_127 : _GEN_7720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_68_T_3 = _myNewVec_127_T_1 + 16'h3b; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_7723 = 7'h1 == _myNewVec_68_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7724 = 7'h2 == _myNewVec_68_T_3[6:0] ? myVec_2 : _GEN_7723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7725 = 7'h3 == _myNewVec_68_T_3[6:0] ? myVec_3 : _GEN_7724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7726 = 7'h4 == _myNewVec_68_T_3[6:0] ? myVec_4 : _GEN_7725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7727 = 7'h5 == _myNewVec_68_T_3[6:0] ? myVec_5 : _GEN_7726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7728 = 7'h6 == _myNewVec_68_T_3[6:0] ? myVec_6 : _GEN_7727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7729 = 7'h7 == _myNewVec_68_T_3[6:0] ? myVec_7 : _GEN_7728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7730 = 7'h8 == _myNewVec_68_T_3[6:0] ? myVec_8 : _GEN_7729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7731 = 7'h9 == _myNewVec_68_T_3[6:0] ? myVec_9 : _GEN_7730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7732 = 7'ha == _myNewVec_68_T_3[6:0] ? myVec_10 : _GEN_7731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7733 = 7'hb == _myNewVec_68_T_3[6:0] ? myVec_11 : _GEN_7732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7734 = 7'hc == _myNewVec_68_T_3[6:0] ? myVec_12 : _GEN_7733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7735 = 7'hd == _myNewVec_68_T_3[6:0] ? myVec_13 : _GEN_7734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7736 = 7'he == _myNewVec_68_T_3[6:0] ? myVec_14 : _GEN_7735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7737 = 7'hf == _myNewVec_68_T_3[6:0] ? myVec_15 : _GEN_7736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7738 = 7'h10 == _myNewVec_68_T_3[6:0] ? myVec_16 : _GEN_7737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7739 = 7'h11 == _myNewVec_68_T_3[6:0] ? myVec_17 : _GEN_7738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7740 = 7'h12 == _myNewVec_68_T_3[6:0] ? myVec_18 : _GEN_7739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7741 = 7'h13 == _myNewVec_68_T_3[6:0] ? myVec_19 : _GEN_7740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7742 = 7'h14 == _myNewVec_68_T_3[6:0] ? myVec_20 : _GEN_7741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7743 = 7'h15 == _myNewVec_68_T_3[6:0] ? myVec_21 : _GEN_7742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7744 = 7'h16 == _myNewVec_68_T_3[6:0] ? myVec_22 : _GEN_7743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7745 = 7'h17 == _myNewVec_68_T_3[6:0] ? myVec_23 : _GEN_7744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7746 = 7'h18 == _myNewVec_68_T_3[6:0] ? myVec_24 : _GEN_7745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7747 = 7'h19 == _myNewVec_68_T_3[6:0] ? myVec_25 : _GEN_7746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7748 = 7'h1a == _myNewVec_68_T_3[6:0] ? myVec_26 : _GEN_7747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7749 = 7'h1b == _myNewVec_68_T_3[6:0] ? myVec_27 : _GEN_7748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7750 = 7'h1c == _myNewVec_68_T_3[6:0] ? myVec_28 : _GEN_7749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7751 = 7'h1d == _myNewVec_68_T_3[6:0] ? myVec_29 : _GEN_7750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7752 = 7'h1e == _myNewVec_68_T_3[6:0] ? myVec_30 : _GEN_7751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7753 = 7'h1f == _myNewVec_68_T_3[6:0] ? myVec_31 : _GEN_7752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7754 = 7'h20 == _myNewVec_68_T_3[6:0] ? myVec_32 : _GEN_7753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7755 = 7'h21 == _myNewVec_68_T_3[6:0] ? myVec_33 : _GEN_7754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7756 = 7'h22 == _myNewVec_68_T_3[6:0] ? myVec_34 : _GEN_7755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7757 = 7'h23 == _myNewVec_68_T_3[6:0] ? myVec_35 : _GEN_7756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7758 = 7'h24 == _myNewVec_68_T_3[6:0] ? myVec_36 : _GEN_7757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7759 = 7'h25 == _myNewVec_68_T_3[6:0] ? myVec_37 : _GEN_7758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7760 = 7'h26 == _myNewVec_68_T_3[6:0] ? myVec_38 : _GEN_7759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7761 = 7'h27 == _myNewVec_68_T_3[6:0] ? myVec_39 : _GEN_7760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7762 = 7'h28 == _myNewVec_68_T_3[6:0] ? myVec_40 : _GEN_7761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7763 = 7'h29 == _myNewVec_68_T_3[6:0] ? myVec_41 : _GEN_7762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7764 = 7'h2a == _myNewVec_68_T_3[6:0] ? myVec_42 : _GEN_7763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7765 = 7'h2b == _myNewVec_68_T_3[6:0] ? myVec_43 : _GEN_7764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7766 = 7'h2c == _myNewVec_68_T_3[6:0] ? myVec_44 : _GEN_7765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7767 = 7'h2d == _myNewVec_68_T_3[6:0] ? myVec_45 : _GEN_7766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7768 = 7'h2e == _myNewVec_68_T_3[6:0] ? myVec_46 : _GEN_7767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7769 = 7'h2f == _myNewVec_68_T_3[6:0] ? myVec_47 : _GEN_7768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7770 = 7'h30 == _myNewVec_68_T_3[6:0] ? myVec_48 : _GEN_7769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7771 = 7'h31 == _myNewVec_68_T_3[6:0] ? myVec_49 : _GEN_7770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7772 = 7'h32 == _myNewVec_68_T_3[6:0] ? myVec_50 : _GEN_7771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7773 = 7'h33 == _myNewVec_68_T_3[6:0] ? myVec_51 : _GEN_7772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7774 = 7'h34 == _myNewVec_68_T_3[6:0] ? myVec_52 : _GEN_7773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7775 = 7'h35 == _myNewVec_68_T_3[6:0] ? myVec_53 : _GEN_7774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7776 = 7'h36 == _myNewVec_68_T_3[6:0] ? myVec_54 : _GEN_7775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7777 = 7'h37 == _myNewVec_68_T_3[6:0] ? myVec_55 : _GEN_7776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7778 = 7'h38 == _myNewVec_68_T_3[6:0] ? myVec_56 : _GEN_7777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7779 = 7'h39 == _myNewVec_68_T_3[6:0] ? myVec_57 : _GEN_7778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7780 = 7'h3a == _myNewVec_68_T_3[6:0] ? myVec_58 : _GEN_7779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7781 = 7'h3b == _myNewVec_68_T_3[6:0] ? myVec_59 : _GEN_7780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7782 = 7'h3c == _myNewVec_68_T_3[6:0] ? myVec_60 : _GEN_7781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7783 = 7'h3d == _myNewVec_68_T_3[6:0] ? myVec_61 : _GEN_7782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7784 = 7'h3e == _myNewVec_68_T_3[6:0] ? myVec_62 : _GEN_7783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7785 = 7'h3f == _myNewVec_68_T_3[6:0] ? myVec_63 : _GEN_7784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7786 = 7'h40 == _myNewVec_68_T_3[6:0] ? myVec_64 : _GEN_7785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7787 = 7'h41 == _myNewVec_68_T_3[6:0] ? myVec_65 : _GEN_7786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7788 = 7'h42 == _myNewVec_68_T_3[6:0] ? myVec_66 : _GEN_7787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7789 = 7'h43 == _myNewVec_68_T_3[6:0] ? myVec_67 : _GEN_7788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7790 = 7'h44 == _myNewVec_68_T_3[6:0] ? myVec_68 : _GEN_7789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7791 = 7'h45 == _myNewVec_68_T_3[6:0] ? myVec_69 : _GEN_7790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7792 = 7'h46 == _myNewVec_68_T_3[6:0] ? myVec_70 : _GEN_7791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7793 = 7'h47 == _myNewVec_68_T_3[6:0] ? myVec_71 : _GEN_7792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7794 = 7'h48 == _myNewVec_68_T_3[6:0] ? myVec_72 : _GEN_7793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7795 = 7'h49 == _myNewVec_68_T_3[6:0] ? myVec_73 : _GEN_7794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7796 = 7'h4a == _myNewVec_68_T_3[6:0] ? myVec_74 : _GEN_7795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7797 = 7'h4b == _myNewVec_68_T_3[6:0] ? myVec_75 : _GEN_7796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7798 = 7'h4c == _myNewVec_68_T_3[6:0] ? myVec_76 : _GEN_7797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7799 = 7'h4d == _myNewVec_68_T_3[6:0] ? myVec_77 : _GEN_7798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7800 = 7'h4e == _myNewVec_68_T_3[6:0] ? myVec_78 : _GEN_7799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7801 = 7'h4f == _myNewVec_68_T_3[6:0] ? myVec_79 : _GEN_7800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7802 = 7'h50 == _myNewVec_68_T_3[6:0] ? myVec_80 : _GEN_7801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7803 = 7'h51 == _myNewVec_68_T_3[6:0] ? myVec_81 : _GEN_7802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7804 = 7'h52 == _myNewVec_68_T_3[6:0] ? myVec_82 : _GEN_7803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7805 = 7'h53 == _myNewVec_68_T_3[6:0] ? myVec_83 : _GEN_7804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7806 = 7'h54 == _myNewVec_68_T_3[6:0] ? myVec_84 : _GEN_7805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7807 = 7'h55 == _myNewVec_68_T_3[6:0] ? myVec_85 : _GEN_7806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7808 = 7'h56 == _myNewVec_68_T_3[6:0] ? myVec_86 : _GEN_7807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7809 = 7'h57 == _myNewVec_68_T_3[6:0] ? myVec_87 : _GEN_7808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7810 = 7'h58 == _myNewVec_68_T_3[6:0] ? myVec_88 : _GEN_7809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7811 = 7'h59 == _myNewVec_68_T_3[6:0] ? myVec_89 : _GEN_7810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7812 = 7'h5a == _myNewVec_68_T_3[6:0] ? myVec_90 : _GEN_7811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7813 = 7'h5b == _myNewVec_68_T_3[6:0] ? myVec_91 : _GEN_7812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7814 = 7'h5c == _myNewVec_68_T_3[6:0] ? myVec_92 : _GEN_7813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7815 = 7'h5d == _myNewVec_68_T_3[6:0] ? myVec_93 : _GEN_7814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7816 = 7'h5e == _myNewVec_68_T_3[6:0] ? myVec_94 : _GEN_7815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7817 = 7'h5f == _myNewVec_68_T_3[6:0] ? myVec_95 : _GEN_7816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7818 = 7'h60 == _myNewVec_68_T_3[6:0] ? myVec_96 : _GEN_7817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7819 = 7'h61 == _myNewVec_68_T_3[6:0] ? myVec_97 : _GEN_7818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7820 = 7'h62 == _myNewVec_68_T_3[6:0] ? myVec_98 : _GEN_7819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7821 = 7'h63 == _myNewVec_68_T_3[6:0] ? myVec_99 : _GEN_7820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7822 = 7'h64 == _myNewVec_68_T_3[6:0] ? myVec_100 : _GEN_7821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7823 = 7'h65 == _myNewVec_68_T_3[6:0] ? myVec_101 : _GEN_7822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7824 = 7'h66 == _myNewVec_68_T_3[6:0] ? myVec_102 : _GEN_7823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7825 = 7'h67 == _myNewVec_68_T_3[6:0] ? myVec_103 : _GEN_7824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7826 = 7'h68 == _myNewVec_68_T_3[6:0] ? myVec_104 : _GEN_7825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7827 = 7'h69 == _myNewVec_68_T_3[6:0] ? myVec_105 : _GEN_7826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7828 = 7'h6a == _myNewVec_68_T_3[6:0] ? myVec_106 : _GEN_7827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7829 = 7'h6b == _myNewVec_68_T_3[6:0] ? myVec_107 : _GEN_7828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7830 = 7'h6c == _myNewVec_68_T_3[6:0] ? myVec_108 : _GEN_7829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7831 = 7'h6d == _myNewVec_68_T_3[6:0] ? myVec_109 : _GEN_7830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7832 = 7'h6e == _myNewVec_68_T_3[6:0] ? myVec_110 : _GEN_7831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7833 = 7'h6f == _myNewVec_68_T_3[6:0] ? myVec_111 : _GEN_7832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7834 = 7'h70 == _myNewVec_68_T_3[6:0] ? myVec_112 : _GEN_7833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7835 = 7'h71 == _myNewVec_68_T_3[6:0] ? myVec_113 : _GEN_7834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7836 = 7'h72 == _myNewVec_68_T_3[6:0] ? myVec_114 : _GEN_7835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7837 = 7'h73 == _myNewVec_68_T_3[6:0] ? myVec_115 : _GEN_7836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7838 = 7'h74 == _myNewVec_68_T_3[6:0] ? myVec_116 : _GEN_7837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7839 = 7'h75 == _myNewVec_68_T_3[6:0] ? myVec_117 : _GEN_7838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7840 = 7'h76 == _myNewVec_68_T_3[6:0] ? myVec_118 : _GEN_7839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7841 = 7'h77 == _myNewVec_68_T_3[6:0] ? myVec_119 : _GEN_7840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7842 = 7'h78 == _myNewVec_68_T_3[6:0] ? myVec_120 : _GEN_7841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7843 = 7'h79 == _myNewVec_68_T_3[6:0] ? myVec_121 : _GEN_7842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7844 = 7'h7a == _myNewVec_68_T_3[6:0] ? myVec_122 : _GEN_7843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7845 = 7'h7b == _myNewVec_68_T_3[6:0] ? myVec_123 : _GEN_7844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7846 = 7'h7c == _myNewVec_68_T_3[6:0] ? myVec_124 : _GEN_7845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7847 = 7'h7d == _myNewVec_68_T_3[6:0] ? myVec_125 : _GEN_7846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7848 = 7'h7e == _myNewVec_68_T_3[6:0] ? myVec_126 : _GEN_7847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_68 = 7'h7f == _myNewVec_68_T_3[6:0] ? myVec_127 : _GEN_7848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_67_T_3 = _myNewVec_127_T_1 + 16'h3c; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_7851 = 7'h1 == _myNewVec_67_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7852 = 7'h2 == _myNewVec_67_T_3[6:0] ? myVec_2 : _GEN_7851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7853 = 7'h3 == _myNewVec_67_T_3[6:0] ? myVec_3 : _GEN_7852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7854 = 7'h4 == _myNewVec_67_T_3[6:0] ? myVec_4 : _GEN_7853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7855 = 7'h5 == _myNewVec_67_T_3[6:0] ? myVec_5 : _GEN_7854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7856 = 7'h6 == _myNewVec_67_T_3[6:0] ? myVec_6 : _GEN_7855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7857 = 7'h7 == _myNewVec_67_T_3[6:0] ? myVec_7 : _GEN_7856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7858 = 7'h8 == _myNewVec_67_T_3[6:0] ? myVec_8 : _GEN_7857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7859 = 7'h9 == _myNewVec_67_T_3[6:0] ? myVec_9 : _GEN_7858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7860 = 7'ha == _myNewVec_67_T_3[6:0] ? myVec_10 : _GEN_7859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7861 = 7'hb == _myNewVec_67_T_3[6:0] ? myVec_11 : _GEN_7860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7862 = 7'hc == _myNewVec_67_T_3[6:0] ? myVec_12 : _GEN_7861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7863 = 7'hd == _myNewVec_67_T_3[6:0] ? myVec_13 : _GEN_7862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7864 = 7'he == _myNewVec_67_T_3[6:0] ? myVec_14 : _GEN_7863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7865 = 7'hf == _myNewVec_67_T_3[6:0] ? myVec_15 : _GEN_7864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7866 = 7'h10 == _myNewVec_67_T_3[6:0] ? myVec_16 : _GEN_7865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7867 = 7'h11 == _myNewVec_67_T_3[6:0] ? myVec_17 : _GEN_7866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7868 = 7'h12 == _myNewVec_67_T_3[6:0] ? myVec_18 : _GEN_7867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7869 = 7'h13 == _myNewVec_67_T_3[6:0] ? myVec_19 : _GEN_7868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7870 = 7'h14 == _myNewVec_67_T_3[6:0] ? myVec_20 : _GEN_7869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7871 = 7'h15 == _myNewVec_67_T_3[6:0] ? myVec_21 : _GEN_7870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7872 = 7'h16 == _myNewVec_67_T_3[6:0] ? myVec_22 : _GEN_7871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7873 = 7'h17 == _myNewVec_67_T_3[6:0] ? myVec_23 : _GEN_7872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7874 = 7'h18 == _myNewVec_67_T_3[6:0] ? myVec_24 : _GEN_7873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7875 = 7'h19 == _myNewVec_67_T_3[6:0] ? myVec_25 : _GEN_7874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7876 = 7'h1a == _myNewVec_67_T_3[6:0] ? myVec_26 : _GEN_7875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7877 = 7'h1b == _myNewVec_67_T_3[6:0] ? myVec_27 : _GEN_7876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7878 = 7'h1c == _myNewVec_67_T_3[6:0] ? myVec_28 : _GEN_7877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7879 = 7'h1d == _myNewVec_67_T_3[6:0] ? myVec_29 : _GEN_7878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7880 = 7'h1e == _myNewVec_67_T_3[6:0] ? myVec_30 : _GEN_7879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7881 = 7'h1f == _myNewVec_67_T_3[6:0] ? myVec_31 : _GEN_7880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7882 = 7'h20 == _myNewVec_67_T_3[6:0] ? myVec_32 : _GEN_7881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7883 = 7'h21 == _myNewVec_67_T_3[6:0] ? myVec_33 : _GEN_7882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7884 = 7'h22 == _myNewVec_67_T_3[6:0] ? myVec_34 : _GEN_7883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7885 = 7'h23 == _myNewVec_67_T_3[6:0] ? myVec_35 : _GEN_7884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7886 = 7'h24 == _myNewVec_67_T_3[6:0] ? myVec_36 : _GEN_7885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7887 = 7'h25 == _myNewVec_67_T_3[6:0] ? myVec_37 : _GEN_7886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7888 = 7'h26 == _myNewVec_67_T_3[6:0] ? myVec_38 : _GEN_7887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7889 = 7'h27 == _myNewVec_67_T_3[6:0] ? myVec_39 : _GEN_7888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7890 = 7'h28 == _myNewVec_67_T_3[6:0] ? myVec_40 : _GEN_7889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7891 = 7'h29 == _myNewVec_67_T_3[6:0] ? myVec_41 : _GEN_7890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7892 = 7'h2a == _myNewVec_67_T_3[6:0] ? myVec_42 : _GEN_7891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7893 = 7'h2b == _myNewVec_67_T_3[6:0] ? myVec_43 : _GEN_7892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7894 = 7'h2c == _myNewVec_67_T_3[6:0] ? myVec_44 : _GEN_7893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7895 = 7'h2d == _myNewVec_67_T_3[6:0] ? myVec_45 : _GEN_7894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7896 = 7'h2e == _myNewVec_67_T_3[6:0] ? myVec_46 : _GEN_7895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7897 = 7'h2f == _myNewVec_67_T_3[6:0] ? myVec_47 : _GEN_7896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7898 = 7'h30 == _myNewVec_67_T_3[6:0] ? myVec_48 : _GEN_7897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7899 = 7'h31 == _myNewVec_67_T_3[6:0] ? myVec_49 : _GEN_7898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7900 = 7'h32 == _myNewVec_67_T_3[6:0] ? myVec_50 : _GEN_7899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7901 = 7'h33 == _myNewVec_67_T_3[6:0] ? myVec_51 : _GEN_7900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7902 = 7'h34 == _myNewVec_67_T_3[6:0] ? myVec_52 : _GEN_7901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7903 = 7'h35 == _myNewVec_67_T_3[6:0] ? myVec_53 : _GEN_7902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7904 = 7'h36 == _myNewVec_67_T_3[6:0] ? myVec_54 : _GEN_7903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7905 = 7'h37 == _myNewVec_67_T_3[6:0] ? myVec_55 : _GEN_7904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7906 = 7'h38 == _myNewVec_67_T_3[6:0] ? myVec_56 : _GEN_7905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7907 = 7'h39 == _myNewVec_67_T_3[6:0] ? myVec_57 : _GEN_7906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7908 = 7'h3a == _myNewVec_67_T_3[6:0] ? myVec_58 : _GEN_7907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7909 = 7'h3b == _myNewVec_67_T_3[6:0] ? myVec_59 : _GEN_7908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7910 = 7'h3c == _myNewVec_67_T_3[6:0] ? myVec_60 : _GEN_7909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7911 = 7'h3d == _myNewVec_67_T_3[6:0] ? myVec_61 : _GEN_7910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7912 = 7'h3e == _myNewVec_67_T_3[6:0] ? myVec_62 : _GEN_7911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7913 = 7'h3f == _myNewVec_67_T_3[6:0] ? myVec_63 : _GEN_7912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7914 = 7'h40 == _myNewVec_67_T_3[6:0] ? myVec_64 : _GEN_7913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7915 = 7'h41 == _myNewVec_67_T_3[6:0] ? myVec_65 : _GEN_7914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7916 = 7'h42 == _myNewVec_67_T_3[6:0] ? myVec_66 : _GEN_7915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7917 = 7'h43 == _myNewVec_67_T_3[6:0] ? myVec_67 : _GEN_7916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7918 = 7'h44 == _myNewVec_67_T_3[6:0] ? myVec_68 : _GEN_7917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7919 = 7'h45 == _myNewVec_67_T_3[6:0] ? myVec_69 : _GEN_7918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7920 = 7'h46 == _myNewVec_67_T_3[6:0] ? myVec_70 : _GEN_7919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7921 = 7'h47 == _myNewVec_67_T_3[6:0] ? myVec_71 : _GEN_7920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7922 = 7'h48 == _myNewVec_67_T_3[6:0] ? myVec_72 : _GEN_7921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7923 = 7'h49 == _myNewVec_67_T_3[6:0] ? myVec_73 : _GEN_7922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7924 = 7'h4a == _myNewVec_67_T_3[6:0] ? myVec_74 : _GEN_7923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7925 = 7'h4b == _myNewVec_67_T_3[6:0] ? myVec_75 : _GEN_7924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7926 = 7'h4c == _myNewVec_67_T_3[6:0] ? myVec_76 : _GEN_7925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7927 = 7'h4d == _myNewVec_67_T_3[6:0] ? myVec_77 : _GEN_7926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7928 = 7'h4e == _myNewVec_67_T_3[6:0] ? myVec_78 : _GEN_7927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7929 = 7'h4f == _myNewVec_67_T_3[6:0] ? myVec_79 : _GEN_7928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7930 = 7'h50 == _myNewVec_67_T_3[6:0] ? myVec_80 : _GEN_7929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7931 = 7'h51 == _myNewVec_67_T_3[6:0] ? myVec_81 : _GEN_7930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7932 = 7'h52 == _myNewVec_67_T_3[6:0] ? myVec_82 : _GEN_7931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7933 = 7'h53 == _myNewVec_67_T_3[6:0] ? myVec_83 : _GEN_7932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7934 = 7'h54 == _myNewVec_67_T_3[6:0] ? myVec_84 : _GEN_7933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7935 = 7'h55 == _myNewVec_67_T_3[6:0] ? myVec_85 : _GEN_7934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7936 = 7'h56 == _myNewVec_67_T_3[6:0] ? myVec_86 : _GEN_7935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7937 = 7'h57 == _myNewVec_67_T_3[6:0] ? myVec_87 : _GEN_7936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7938 = 7'h58 == _myNewVec_67_T_3[6:0] ? myVec_88 : _GEN_7937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7939 = 7'h59 == _myNewVec_67_T_3[6:0] ? myVec_89 : _GEN_7938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7940 = 7'h5a == _myNewVec_67_T_3[6:0] ? myVec_90 : _GEN_7939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7941 = 7'h5b == _myNewVec_67_T_3[6:0] ? myVec_91 : _GEN_7940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7942 = 7'h5c == _myNewVec_67_T_3[6:0] ? myVec_92 : _GEN_7941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7943 = 7'h5d == _myNewVec_67_T_3[6:0] ? myVec_93 : _GEN_7942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7944 = 7'h5e == _myNewVec_67_T_3[6:0] ? myVec_94 : _GEN_7943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7945 = 7'h5f == _myNewVec_67_T_3[6:0] ? myVec_95 : _GEN_7944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7946 = 7'h60 == _myNewVec_67_T_3[6:0] ? myVec_96 : _GEN_7945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7947 = 7'h61 == _myNewVec_67_T_3[6:0] ? myVec_97 : _GEN_7946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7948 = 7'h62 == _myNewVec_67_T_3[6:0] ? myVec_98 : _GEN_7947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7949 = 7'h63 == _myNewVec_67_T_3[6:0] ? myVec_99 : _GEN_7948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7950 = 7'h64 == _myNewVec_67_T_3[6:0] ? myVec_100 : _GEN_7949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7951 = 7'h65 == _myNewVec_67_T_3[6:0] ? myVec_101 : _GEN_7950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7952 = 7'h66 == _myNewVec_67_T_3[6:0] ? myVec_102 : _GEN_7951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7953 = 7'h67 == _myNewVec_67_T_3[6:0] ? myVec_103 : _GEN_7952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7954 = 7'h68 == _myNewVec_67_T_3[6:0] ? myVec_104 : _GEN_7953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7955 = 7'h69 == _myNewVec_67_T_3[6:0] ? myVec_105 : _GEN_7954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7956 = 7'h6a == _myNewVec_67_T_3[6:0] ? myVec_106 : _GEN_7955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7957 = 7'h6b == _myNewVec_67_T_3[6:0] ? myVec_107 : _GEN_7956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7958 = 7'h6c == _myNewVec_67_T_3[6:0] ? myVec_108 : _GEN_7957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7959 = 7'h6d == _myNewVec_67_T_3[6:0] ? myVec_109 : _GEN_7958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7960 = 7'h6e == _myNewVec_67_T_3[6:0] ? myVec_110 : _GEN_7959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7961 = 7'h6f == _myNewVec_67_T_3[6:0] ? myVec_111 : _GEN_7960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7962 = 7'h70 == _myNewVec_67_T_3[6:0] ? myVec_112 : _GEN_7961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7963 = 7'h71 == _myNewVec_67_T_3[6:0] ? myVec_113 : _GEN_7962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7964 = 7'h72 == _myNewVec_67_T_3[6:0] ? myVec_114 : _GEN_7963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7965 = 7'h73 == _myNewVec_67_T_3[6:0] ? myVec_115 : _GEN_7964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7966 = 7'h74 == _myNewVec_67_T_3[6:0] ? myVec_116 : _GEN_7965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7967 = 7'h75 == _myNewVec_67_T_3[6:0] ? myVec_117 : _GEN_7966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7968 = 7'h76 == _myNewVec_67_T_3[6:0] ? myVec_118 : _GEN_7967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7969 = 7'h77 == _myNewVec_67_T_3[6:0] ? myVec_119 : _GEN_7968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7970 = 7'h78 == _myNewVec_67_T_3[6:0] ? myVec_120 : _GEN_7969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7971 = 7'h79 == _myNewVec_67_T_3[6:0] ? myVec_121 : _GEN_7970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7972 = 7'h7a == _myNewVec_67_T_3[6:0] ? myVec_122 : _GEN_7971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7973 = 7'h7b == _myNewVec_67_T_3[6:0] ? myVec_123 : _GEN_7972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7974 = 7'h7c == _myNewVec_67_T_3[6:0] ? myVec_124 : _GEN_7973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7975 = 7'h7d == _myNewVec_67_T_3[6:0] ? myVec_125 : _GEN_7974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7976 = 7'h7e == _myNewVec_67_T_3[6:0] ? myVec_126 : _GEN_7975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_67 = 7'h7f == _myNewVec_67_T_3[6:0] ? myVec_127 : _GEN_7976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_66_T_3 = _myNewVec_127_T_1 + 16'h3d; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_7979 = 7'h1 == _myNewVec_66_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7980 = 7'h2 == _myNewVec_66_T_3[6:0] ? myVec_2 : _GEN_7979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7981 = 7'h3 == _myNewVec_66_T_3[6:0] ? myVec_3 : _GEN_7980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7982 = 7'h4 == _myNewVec_66_T_3[6:0] ? myVec_4 : _GEN_7981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7983 = 7'h5 == _myNewVec_66_T_3[6:0] ? myVec_5 : _GEN_7982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7984 = 7'h6 == _myNewVec_66_T_3[6:0] ? myVec_6 : _GEN_7983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7985 = 7'h7 == _myNewVec_66_T_3[6:0] ? myVec_7 : _GEN_7984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7986 = 7'h8 == _myNewVec_66_T_3[6:0] ? myVec_8 : _GEN_7985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7987 = 7'h9 == _myNewVec_66_T_3[6:0] ? myVec_9 : _GEN_7986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7988 = 7'ha == _myNewVec_66_T_3[6:0] ? myVec_10 : _GEN_7987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7989 = 7'hb == _myNewVec_66_T_3[6:0] ? myVec_11 : _GEN_7988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7990 = 7'hc == _myNewVec_66_T_3[6:0] ? myVec_12 : _GEN_7989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7991 = 7'hd == _myNewVec_66_T_3[6:0] ? myVec_13 : _GEN_7990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7992 = 7'he == _myNewVec_66_T_3[6:0] ? myVec_14 : _GEN_7991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7993 = 7'hf == _myNewVec_66_T_3[6:0] ? myVec_15 : _GEN_7992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7994 = 7'h10 == _myNewVec_66_T_3[6:0] ? myVec_16 : _GEN_7993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7995 = 7'h11 == _myNewVec_66_T_3[6:0] ? myVec_17 : _GEN_7994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7996 = 7'h12 == _myNewVec_66_T_3[6:0] ? myVec_18 : _GEN_7995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7997 = 7'h13 == _myNewVec_66_T_3[6:0] ? myVec_19 : _GEN_7996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7998 = 7'h14 == _myNewVec_66_T_3[6:0] ? myVec_20 : _GEN_7997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_7999 = 7'h15 == _myNewVec_66_T_3[6:0] ? myVec_21 : _GEN_7998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8000 = 7'h16 == _myNewVec_66_T_3[6:0] ? myVec_22 : _GEN_7999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8001 = 7'h17 == _myNewVec_66_T_3[6:0] ? myVec_23 : _GEN_8000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8002 = 7'h18 == _myNewVec_66_T_3[6:0] ? myVec_24 : _GEN_8001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8003 = 7'h19 == _myNewVec_66_T_3[6:0] ? myVec_25 : _GEN_8002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8004 = 7'h1a == _myNewVec_66_T_3[6:0] ? myVec_26 : _GEN_8003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8005 = 7'h1b == _myNewVec_66_T_3[6:0] ? myVec_27 : _GEN_8004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8006 = 7'h1c == _myNewVec_66_T_3[6:0] ? myVec_28 : _GEN_8005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8007 = 7'h1d == _myNewVec_66_T_3[6:0] ? myVec_29 : _GEN_8006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8008 = 7'h1e == _myNewVec_66_T_3[6:0] ? myVec_30 : _GEN_8007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8009 = 7'h1f == _myNewVec_66_T_3[6:0] ? myVec_31 : _GEN_8008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8010 = 7'h20 == _myNewVec_66_T_3[6:0] ? myVec_32 : _GEN_8009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8011 = 7'h21 == _myNewVec_66_T_3[6:0] ? myVec_33 : _GEN_8010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8012 = 7'h22 == _myNewVec_66_T_3[6:0] ? myVec_34 : _GEN_8011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8013 = 7'h23 == _myNewVec_66_T_3[6:0] ? myVec_35 : _GEN_8012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8014 = 7'h24 == _myNewVec_66_T_3[6:0] ? myVec_36 : _GEN_8013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8015 = 7'h25 == _myNewVec_66_T_3[6:0] ? myVec_37 : _GEN_8014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8016 = 7'h26 == _myNewVec_66_T_3[6:0] ? myVec_38 : _GEN_8015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8017 = 7'h27 == _myNewVec_66_T_3[6:0] ? myVec_39 : _GEN_8016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8018 = 7'h28 == _myNewVec_66_T_3[6:0] ? myVec_40 : _GEN_8017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8019 = 7'h29 == _myNewVec_66_T_3[6:0] ? myVec_41 : _GEN_8018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8020 = 7'h2a == _myNewVec_66_T_3[6:0] ? myVec_42 : _GEN_8019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8021 = 7'h2b == _myNewVec_66_T_3[6:0] ? myVec_43 : _GEN_8020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8022 = 7'h2c == _myNewVec_66_T_3[6:0] ? myVec_44 : _GEN_8021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8023 = 7'h2d == _myNewVec_66_T_3[6:0] ? myVec_45 : _GEN_8022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8024 = 7'h2e == _myNewVec_66_T_3[6:0] ? myVec_46 : _GEN_8023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8025 = 7'h2f == _myNewVec_66_T_3[6:0] ? myVec_47 : _GEN_8024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8026 = 7'h30 == _myNewVec_66_T_3[6:0] ? myVec_48 : _GEN_8025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8027 = 7'h31 == _myNewVec_66_T_3[6:0] ? myVec_49 : _GEN_8026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8028 = 7'h32 == _myNewVec_66_T_3[6:0] ? myVec_50 : _GEN_8027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8029 = 7'h33 == _myNewVec_66_T_3[6:0] ? myVec_51 : _GEN_8028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8030 = 7'h34 == _myNewVec_66_T_3[6:0] ? myVec_52 : _GEN_8029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8031 = 7'h35 == _myNewVec_66_T_3[6:0] ? myVec_53 : _GEN_8030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8032 = 7'h36 == _myNewVec_66_T_3[6:0] ? myVec_54 : _GEN_8031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8033 = 7'h37 == _myNewVec_66_T_3[6:0] ? myVec_55 : _GEN_8032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8034 = 7'h38 == _myNewVec_66_T_3[6:0] ? myVec_56 : _GEN_8033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8035 = 7'h39 == _myNewVec_66_T_3[6:0] ? myVec_57 : _GEN_8034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8036 = 7'h3a == _myNewVec_66_T_3[6:0] ? myVec_58 : _GEN_8035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8037 = 7'h3b == _myNewVec_66_T_3[6:0] ? myVec_59 : _GEN_8036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8038 = 7'h3c == _myNewVec_66_T_3[6:0] ? myVec_60 : _GEN_8037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8039 = 7'h3d == _myNewVec_66_T_3[6:0] ? myVec_61 : _GEN_8038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8040 = 7'h3e == _myNewVec_66_T_3[6:0] ? myVec_62 : _GEN_8039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8041 = 7'h3f == _myNewVec_66_T_3[6:0] ? myVec_63 : _GEN_8040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8042 = 7'h40 == _myNewVec_66_T_3[6:0] ? myVec_64 : _GEN_8041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8043 = 7'h41 == _myNewVec_66_T_3[6:0] ? myVec_65 : _GEN_8042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8044 = 7'h42 == _myNewVec_66_T_3[6:0] ? myVec_66 : _GEN_8043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8045 = 7'h43 == _myNewVec_66_T_3[6:0] ? myVec_67 : _GEN_8044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8046 = 7'h44 == _myNewVec_66_T_3[6:0] ? myVec_68 : _GEN_8045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8047 = 7'h45 == _myNewVec_66_T_3[6:0] ? myVec_69 : _GEN_8046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8048 = 7'h46 == _myNewVec_66_T_3[6:0] ? myVec_70 : _GEN_8047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8049 = 7'h47 == _myNewVec_66_T_3[6:0] ? myVec_71 : _GEN_8048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8050 = 7'h48 == _myNewVec_66_T_3[6:0] ? myVec_72 : _GEN_8049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8051 = 7'h49 == _myNewVec_66_T_3[6:0] ? myVec_73 : _GEN_8050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8052 = 7'h4a == _myNewVec_66_T_3[6:0] ? myVec_74 : _GEN_8051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8053 = 7'h4b == _myNewVec_66_T_3[6:0] ? myVec_75 : _GEN_8052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8054 = 7'h4c == _myNewVec_66_T_3[6:0] ? myVec_76 : _GEN_8053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8055 = 7'h4d == _myNewVec_66_T_3[6:0] ? myVec_77 : _GEN_8054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8056 = 7'h4e == _myNewVec_66_T_3[6:0] ? myVec_78 : _GEN_8055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8057 = 7'h4f == _myNewVec_66_T_3[6:0] ? myVec_79 : _GEN_8056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8058 = 7'h50 == _myNewVec_66_T_3[6:0] ? myVec_80 : _GEN_8057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8059 = 7'h51 == _myNewVec_66_T_3[6:0] ? myVec_81 : _GEN_8058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8060 = 7'h52 == _myNewVec_66_T_3[6:0] ? myVec_82 : _GEN_8059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8061 = 7'h53 == _myNewVec_66_T_3[6:0] ? myVec_83 : _GEN_8060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8062 = 7'h54 == _myNewVec_66_T_3[6:0] ? myVec_84 : _GEN_8061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8063 = 7'h55 == _myNewVec_66_T_3[6:0] ? myVec_85 : _GEN_8062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8064 = 7'h56 == _myNewVec_66_T_3[6:0] ? myVec_86 : _GEN_8063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8065 = 7'h57 == _myNewVec_66_T_3[6:0] ? myVec_87 : _GEN_8064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8066 = 7'h58 == _myNewVec_66_T_3[6:0] ? myVec_88 : _GEN_8065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8067 = 7'h59 == _myNewVec_66_T_3[6:0] ? myVec_89 : _GEN_8066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8068 = 7'h5a == _myNewVec_66_T_3[6:0] ? myVec_90 : _GEN_8067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8069 = 7'h5b == _myNewVec_66_T_3[6:0] ? myVec_91 : _GEN_8068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8070 = 7'h5c == _myNewVec_66_T_3[6:0] ? myVec_92 : _GEN_8069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8071 = 7'h5d == _myNewVec_66_T_3[6:0] ? myVec_93 : _GEN_8070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8072 = 7'h5e == _myNewVec_66_T_3[6:0] ? myVec_94 : _GEN_8071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8073 = 7'h5f == _myNewVec_66_T_3[6:0] ? myVec_95 : _GEN_8072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8074 = 7'h60 == _myNewVec_66_T_3[6:0] ? myVec_96 : _GEN_8073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8075 = 7'h61 == _myNewVec_66_T_3[6:0] ? myVec_97 : _GEN_8074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8076 = 7'h62 == _myNewVec_66_T_3[6:0] ? myVec_98 : _GEN_8075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8077 = 7'h63 == _myNewVec_66_T_3[6:0] ? myVec_99 : _GEN_8076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8078 = 7'h64 == _myNewVec_66_T_3[6:0] ? myVec_100 : _GEN_8077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8079 = 7'h65 == _myNewVec_66_T_3[6:0] ? myVec_101 : _GEN_8078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8080 = 7'h66 == _myNewVec_66_T_3[6:0] ? myVec_102 : _GEN_8079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8081 = 7'h67 == _myNewVec_66_T_3[6:0] ? myVec_103 : _GEN_8080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8082 = 7'h68 == _myNewVec_66_T_3[6:0] ? myVec_104 : _GEN_8081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8083 = 7'h69 == _myNewVec_66_T_3[6:0] ? myVec_105 : _GEN_8082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8084 = 7'h6a == _myNewVec_66_T_3[6:0] ? myVec_106 : _GEN_8083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8085 = 7'h6b == _myNewVec_66_T_3[6:0] ? myVec_107 : _GEN_8084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8086 = 7'h6c == _myNewVec_66_T_3[6:0] ? myVec_108 : _GEN_8085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8087 = 7'h6d == _myNewVec_66_T_3[6:0] ? myVec_109 : _GEN_8086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8088 = 7'h6e == _myNewVec_66_T_3[6:0] ? myVec_110 : _GEN_8087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8089 = 7'h6f == _myNewVec_66_T_3[6:0] ? myVec_111 : _GEN_8088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8090 = 7'h70 == _myNewVec_66_T_3[6:0] ? myVec_112 : _GEN_8089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8091 = 7'h71 == _myNewVec_66_T_3[6:0] ? myVec_113 : _GEN_8090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8092 = 7'h72 == _myNewVec_66_T_3[6:0] ? myVec_114 : _GEN_8091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8093 = 7'h73 == _myNewVec_66_T_3[6:0] ? myVec_115 : _GEN_8092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8094 = 7'h74 == _myNewVec_66_T_3[6:0] ? myVec_116 : _GEN_8093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8095 = 7'h75 == _myNewVec_66_T_3[6:0] ? myVec_117 : _GEN_8094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8096 = 7'h76 == _myNewVec_66_T_3[6:0] ? myVec_118 : _GEN_8095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8097 = 7'h77 == _myNewVec_66_T_3[6:0] ? myVec_119 : _GEN_8096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8098 = 7'h78 == _myNewVec_66_T_3[6:0] ? myVec_120 : _GEN_8097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8099 = 7'h79 == _myNewVec_66_T_3[6:0] ? myVec_121 : _GEN_8098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8100 = 7'h7a == _myNewVec_66_T_3[6:0] ? myVec_122 : _GEN_8099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8101 = 7'h7b == _myNewVec_66_T_3[6:0] ? myVec_123 : _GEN_8100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8102 = 7'h7c == _myNewVec_66_T_3[6:0] ? myVec_124 : _GEN_8101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8103 = 7'h7d == _myNewVec_66_T_3[6:0] ? myVec_125 : _GEN_8102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8104 = 7'h7e == _myNewVec_66_T_3[6:0] ? myVec_126 : _GEN_8103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_66 = 7'h7f == _myNewVec_66_T_3[6:0] ? myVec_127 : _GEN_8104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_65_T_3 = _myNewVec_127_T_1 + 16'h3e; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_8107 = 7'h1 == _myNewVec_65_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8108 = 7'h2 == _myNewVec_65_T_3[6:0] ? myVec_2 : _GEN_8107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8109 = 7'h3 == _myNewVec_65_T_3[6:0] ? myVec_3 : _GEN_8108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8110 = 7'h4 == _myNewVec_65_T_3[6:0] ? myVec_4 : _GEN_8109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8111 = 7'h5 == _myNewVec_65_T_3[6:0] ? myVec_5 : _GEN_8110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8112 = 7'h6 == _myNewVec_65_T_3[6:0] ? myVec_6 : _GEN_8111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8113 = 7'h7 == _myNewVec_65_T_3[6:0] ? myVec_7 : _GEN_8112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8114 = 7'h8 == _myNewVec_65_T_3[6:0] ? myVec_8 : _GEN_8113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8115 = 7'h9 == _myNewVec_65_T_3[6:0] ? myVec_9 : _GEN_8114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8116 = 7'ha == _myNewVec_65_T_3[6:0] ? myVec_10 : _GEN_8115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8117 = 7'hb == _myNewVec_65_T_3[6:0] ? myVec_11 : _GEN_8116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8118 = 7'hc == _myNewVec_65_T_3[6:0] ? myVec_12 : _GEN_8117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8119 = 7'hd == _myNewVec_65_T_3[6:0] ? myVec_13 : _GEN_8118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8120 = 7'he == _myNewVec_65_T_3[6:0] ? myVec_14 : _GEN_8119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8121 = 7'hf == _myNewVec_65_T_3[6:0] ? myVec_15 : _GEN_8120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8122 = 7'h10 == _myNewVec_65_T_3[6:0] ? myVec_16 : _GEN_8121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8123 = 7'h11 == _myNewVec_65_T_3[6:0] ? myVec_17 : _GEN_8122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8124 = 7'h12 == _myNewVec_65_T_3[6:0] ? myVec_18 : _GEN_8123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8125 = 7'h13 == _myNewVec_65_T_3[6:0] ? myVec_19 : _GEN_8124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8126 = 7'h14 == _myNewVec_65_T_3[6:0] ? myVec_20 : _GEN_8125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8127 = 7'h15 == _myNewVec_65_T_3[6:0] ? myVec_21 : _GEN_8126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8128 = 7'h16 == _myNewVec_65_T_3[6:0] ? myVec_22 : _GEN_8127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8129 = 7'h17 == _myNewVec_65_T_3[6:0] ? myVec_23 : _GEN_8128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8130 = 7'h18 == _myNewVec_65_T_3[6:0] ? myVec_24 : _GEN_8129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8131 = 7'h19 == _myNewVec_65_T_3[6:0] ? myVec_25 : _GEN_8130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8132 = 7'h1a == _myNewVec_65_T_3[6:0] ? myVec_26 : _GEN_8131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8133 = 7'h1b == _myNewVec_65_T_3[6:0] ? myVec_27 : _GEN_8132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8134 = 7'h1c == _myNewVec_65_T_3[6:0] ? myVec_28 : _GEN_8133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8135 = 7'h1d == _myNewVec_65_T_3[6:0] ? myVec_29 : _GEN_8134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8136 = 7'h1e == _myNewVec_65_T_3[6:0] ? myVec_30 : _GEN_8135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8137 = 7'h1f == _myNewVec_65_T_3[6:0] ? myVec_31 : _GEN_8136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8138 = 7'h20 == _myNewVec_65_T_3[6:0] ? myVec_32 : _GEN_8137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8139 = 7'h21 == _myNewVec_65_T_3[6:0] ? myVec_33 : _GEN_8138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8140 = 7'h22 == _myNewVec_65_T_3[6:0] ? myVec_34 : _GEN_8139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8141 = 7'h23 == _myNewVec_65_T_3[6:0] ? myVec_35 : _GEN_8140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8142 = 7'h24 == _myNewVec_65_T_3[6:0] ? myVec_36 : _GEN_8141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8143 = 7'h25 == _myNewVec_65_T_3[6:0] ? myVec_37 : _GEN_8142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8144 = 7'h26 == _myNewVec_65_T_3[6:0] ? myVec_38 : _GEN_8143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8145 = 7'h27 == _myNewVec_65_T_3[6:0] ? myVec_39 : _GEN_8144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8146 = 7'h28 == _myNewVec_65_T_3[6:0] ? myVec_40 : _GEN_8145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8147 = 7'h29 == _myNewVec_65_T_3[6:0] ? myVec_41 : _GEN_8146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8148 = 7'h2a == _myNewVec_65_T_3[6:0] ? myVec_42 : _GEN_8147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8149 = 7'h2b == _myNewVec_65_T_3[6:0] ? myVec_43 : _GEN_8148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8150 = 7'h2c == _myNewVec_65_T_3[6:0] ? myVec_44 : _GEN_8149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8151 = 7'h2d == _myNewVec_65_T_3[6:0] ? myVec_45 : _GEN_8150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8152 = 7'h2e == _myNewVec_65_T_3[6:0] ? myVec_46 : _GEN_8151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8153 = 7'h2f == _myNewVec_65_T_3[6:0] ? myVec_47 : _GEN_8152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8154 = 7'h30 == _myNewVec_65_T_3[6:0] ? myVec_48 : _GEN_8153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8155 = 7'h31 == _myNewVec_65_T_3[6:0] ? myVec_49 : _GEN_8154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8156 = 7'h32 == _myNewVec_65_T_3[6:0] ? myVec_50 : _GEN_8155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8157 = 7'h33 == _myNewVec_65_T_3[6:0] ? myVec_51 : _GEN_8156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8158 = 7'h34 == _myNewVec_65_T_3[6:0] ? myVec_52 : _GEN_8157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8159 = 7'h35 == _myNewVec_65_T_3[6:0] ? myVec_53 : _GEN_8158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8160 = 7'h36 == _myNewVec_65_T_3[6:0] ? myVec_54 : _GEN_8159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8161 = 7'h37 == _myNewVec_65_T_3[6:0] ? myVec_55 : _GEN_8160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8162 = 7'h38 == _myNewVec_65_T_3[6:0] ? myVec_56 : _GEN_8161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8163 = 7'h39 == _myNewVec_65_T_3[6:0] ? myVec_57 : _GEN_8162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8164 = 7'h3a == _myNewVec_65_T_3[6:0] ? myVec_58 : _GEN_8163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8165 = 7'h3b == _myNewVec_65_T_3[6:0] ? myVec_59 : _GEN_8164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8166 = 7'h3c == _myNewVec_65_T_3[6:0] ? myVec_60 : _GEN_8165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8167 = 7'h3d == _myNewVec_65_T_3[6:0] ? myVec_61 : _GEN_8166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8168 = 7'h3e == _myNewVec_65_T_3[6:0] ? myVec_62 : _GEN_8167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8169 = 7'h3f == _myNewVec_65_T_3[6:0] ? myVec_63 : _GEN_8168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8170 = 7'h40 == _myNewVec_65_T_3[6:0] ? myVec_64 : _GEN_8169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8171 = 7'h41 == _myNewVec_65_T_3[6:0] ? myVec_65 : _GEN_8170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8172 = 7'h42 == _myNewVec_65_T_3[6:0] ? myVec_66 : _GEN_8171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8173 = 7'h43 == _myNewVec_65_T_3[6:0] ? myVec_67 : _GEN_8172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8174 = 7'h44 == _myNewVec_65_T_3[6:0] ? myVec_68 : _GEN_8173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8175 = 7'h45 == _myNewVec_65_T_3[6:0] ? myVec_69 : _GEN_8174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8176 = 7'h46 == _myNewVec_65_T_3[6:0] ? myVec_70 : _GEN_8175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8177 = 7'h47 == _myNewVec_65_T_3[6:0] ? myVec_71 : _GEN_8176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8178 = 7'h48 == _myNewVec_65_T_3[6:0] ? myVec_72 : _GEN_8177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8179 = 7'h49 == _myNewVec_65_T_3[6:0] ? myVec_73 : _GEN_8178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8180 = 7'h4a == _myNewVec_65_T_3[6:0] ? myVec_74 : _GEN_8179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8181 = 7'h4b == _myNewVec_65_T_3[6:0] ? myVec_75 : _GEN_8180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8182 = 7'h4c == _myNewVec_65_T_3[6:0] ? myVec_76 : _GEN_8181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8183 = 7'h4d == _myNewVec_65_T_3[6:0] ? myVec_77 : _GEN_8182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8184 = 7'h4e == _myNewVec_65_T_3[6:0] ? myVec_78 : _GEN_8183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8185 = 7'h4f == _myNewVec_65_T_3[6:0] ? myVec_79 : _GEN_8184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8186 = 7'h50 == _myNewVec_65_T_3[6:0] ? myVec_80 : _GEN_8185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8187 = 7'h51 == _myNewVec_65_T_3[6:0] ? myVec_81 : _GEN_8186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8188 = 7'h52 == _myNewVec_65_T_3[6:0] ? myVec_82 : _GEN_8187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8189 = 7'h53 == _myNewVec_65_T_3[6:0] ? myVec_83 : _GEN_8188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8190 = 7'h54 == _myNewVec_65_T_3[6:0] ? myVec_84 : _GEN_8189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8191 = 7'h55 == _myNewVec_65_T_3[6:0] ? myVec_85 : _GEN_8190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8192 = 7'h56 == _myNewVec_65_T_3[6:0] ? myVec_86 : _GEN_8191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8193 = 7'h57 == _myNewVec_65_T_3[6:0] ? myVec_87 : _GEN_8192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8194 = 7'h58 == _myNewVec_65_T_3[6:0] ? myVec_88 : _GEN_8193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8195 = 7'h59 == _myNewVec_65_T_3[6:0] ? myVec_89 : _GEN_8194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8196 = 7'h5a == _myNewVec_65_T_3[6:0] ? myVec_90 : _GEN_8195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8197 = 7'h5b == _myNewVec_65_T_3[6:0] ? myVec_91 : _GEN_8196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8198 = 7'h5c == _myNewVec_65_T_3[6:0] ? myVec_92 : _GEN_8197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8199 = 7'h5d == _myNewVec_65_T_3[6:0] ? myVec_93 : _GEN_8198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8200 = 7'h5e == _myNewVec_65_T_3[6:0] ? myVec_94 : _GEN_8199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8201 = 7'h5f == _myNewVec_65_T_3[6:0] ? myVec_95 : _GEN_8200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8202 = 7'h60 == _myNewVec_65_T_3[6:0] ? myVec_96 : _GEN_8201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8203 = 7'h61 == _myNewVec_65_T_3[6:0] ? myVec_97 : _GEN_8202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8204 = 7'h62 == _myNewVec_65_T_3[6:0] ? myVec_98 : _GEN_8203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8205 = 7'h63 == _myNewVec_65_T_3[6:0] ? myVec_99 : _GEN_8204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8206 = 7'h64 == _myNewVec_65_T_3[6:0] ? myVec_100 : _GEN_8205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8207 = 7'h65 == _myNewVec_65_T_3[6:0] ? myVec_101 : _GEN_8206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8208 = 7'h66 == _myNewVec_65_T_3[6:0] ? myVec_102 : _GEN_8207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8209 = 7'h67 == _myNewVec_65_T_3[6:0] ? myVec_103 : _GEN_8208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8210 = 7'h68 == _myNewVec_65_T_3[6:0] ? myVec_104 : _GEN_8209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8211 = 7'h69 == _myNewVec_65_T_3[6:0] ? myVec_105 : _GEN_8210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8212 = 7'h6a == _myNewVec_65_T_3[6:0] ? myVec_106 : _GEN_8211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8213 = 7'h6b == _myNewVec_65_T_3[6:0] ? myVec_107 : _GEN_8212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8214 = 7'h6c == _myNewVec_65_T_3[6:0] ? myVec_108 : _GEN_8213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8215 = 7'h6d == _myNewVec_65_T_3[6:0] ? myVec_109 : _GEN_8214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8216 = 7'h6e == _myNewVec_65_T_3[6:0] ? myVec_110 : _GEN_8215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8217 = 7'h6f == _myNewVec_65_T_3[6:0] ? myVec_111 : _GEN_8216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8218 = 7'h70 == _myNewVec_65_T_3[6:0] ? myVec_112 : _GEN_8217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8219 = 7'h71 == _myNewVec_65_T_3[6:0] ? myVec_113 : _GEN_8218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8220 = 7'h72 == _myNewVec_65_T_3[6:0] ? myVec_114 : _GEN_8219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8221 = 7'h73 == _myNewVec_65_T_3[6:0] ? myVec_115 : _GEN_8220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8222 = 7'h74 == _myNewVec_65_T_3[6:0] ? myVec_116 : _GEN_8221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8223 = 7'h75 == _myNewVec_65_T_3[6:0] ? myVec_117 : _GEN_8222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8224 = 7'h76 == _myNewVec_65_T_3[6:0] ? myVec_118 : _GEN_8223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8225 = 7'h77 == _myNewVec_65_T_3[6:0] ? myVec_119 : _GEN_8224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8226 = 7'h78 == _myNewVec_65_T_3[6:0] ? myVec_120 : _GEN_8225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8227 = 7'h79 == _myNewVec_65_T_3[6:0] ? myVec_121 : _GEN_8226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8228 = 7'h7a == _myNewVec_65_T_3[6:0] ? myVec_122 : _GEN_8227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8229 = 7'h7b == _myNewVec_65_T_3[6:0] ? myVec_123 : _GEN_8228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8230 = 7'h7c == _myNewVec_65_T_3[6:0] ? myVec_124 : _GEN_8229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8231 = 7'h7d == _myNewVec_65_T_3[6:0] ? myVec_125 : _GEN_8230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8232 = 7'h7e == _myNewVec_65_T_3[6:0] ? myVec_126 : _GEN_8231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_65 = 7'h7f == _myNewVec_65_T_3[6:0] ? myVec_127 : _GEN_8232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_64_T_3 = _myNewVec_127_T_1 + 16'h3f; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_8235 = 7'h1 == _myNewVec_64_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8236 = 7'h2 == _myNewVec_64_T_3[6:0] ? myVec_2 : _GEN_8235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8237 = 7'h3 == _myNewVec_64_T_3[6:0] ? myVec_3 : _GEN_8236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8238 = 7'h4 == _myNewVec_64_T_3[6:0] ? myVec_4 : _GEN_8237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8239 = 7'h5 == _myNewVec_64_T_3[6:0] ? myVec_5 : _GEN_8238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8240 = 7'h6 == _myNewVec_64_T_3[6:0] ? myVec_6 : _GEN_8239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8241 = 7'h7 == _myNewVec_64_T_3[6:0] ? myVec_7 : _GEN_8240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8242 = 7'h8 == _myNewVec_64_T_3[6:0] ? myVec_8 : _GEN_8241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8243 = 7'h9 == _myNewVec_64_T_3[6:0] ? myVec_9 : _GEN_8242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8244 = 7'ha == _myNewVec_64_T_3[6:0] ? myVec_10 : _GEN_8243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8245 = 7'hb == _myNewVec_64_T_3[6:0] ? myVec_11 : _GEN_8244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8246 = 7'hc == _myNewVec_64_T_3[6:0] ? myVec_12 : _GEN_8245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8247 = 7'hd == _myNewVec_64_T_3[6:0] ? myVec_13 : _GEN_8246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8248 = 7'he == _myNewVec_64_T_3[6:0] ? myVec_14 : _GEN_8247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8249 = 7'hf == _myNewVec_64_T_3[6:0] ? myVec_15 : _GEN_8248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8250 = 7'h10 == _myNewVec_64_T_3[6:0] ? myVec_16 : _GEN_8249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8251 = 7'h11 == _myNewVec_64_T_3[6:0] ? myVec_17 : _GEN_8250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8252 = 7'h12 == _myNewVec_64_T_3[6:0] ? myVec_18 : _GEN_8251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8253 = 7'h13 == _myNewVec_64_T_3[6:0] ? myVec_19 : _GEN_8252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8254 = 7'h14 == _myNewVec_64_T_3[6:0] ? myVec_20 : _GEN_8253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8255 = 7'h15 == _myNewVec_64_T_3[6:0] ? myVec_21 : _GEN_8254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8256 = 7'h16 == _myNewVec_64_T_3[6:0] ? myVec_22 : _GEN_8255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8257 = 7'h17 == _myNewVec_64_T_3[6:0] ? myVec_23 : _GEN_8256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8258 = 7'h18 == _myNewVec_64_T_3[6:0] ? myVec_24 : _GEN_8257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8259 = 7'h19 == _myNewVec_64_T_3[6:0] ? myVec_25 : _GEN_8258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8260 = 7'h1a == _myNewVec_64_T_3[6:0] ? myVec_26 : _GEN_8259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8261 = 7'h1b == _myNewVec_64_T_3[6:0] ? myVec_27 : _GEN_8260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8262 = 7'h1c == _myNewVec_64_T_3[6:0] ? myVec_28 : _GEN_8261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8263 = 7'h1d == _myNewVec_64_T_3[6:0] ? myVec_29 : _GEN_8262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8264 = 7'h1e == _myNewVec_64_T_3[6:0] ? myVec_30 : _GEN_8263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8265 = 7'h1f == _myNewVec_64_T_3[6:0] ? myVec_31 : _GEN_8264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8266 = 7'h20 == _myNewVec_64_T_3[6:0] ? myVec_32 : _GEN_8265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8267 = 7'h21 == _myNewVec_64_T_3[6:0] ? myVec_33 : _GEN_8266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8268 = 7'h22 == _myNewVec_64_T_3[6:0] ? myVec_34 : _GEN_8267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8269 = 7'h23 == _myNewVec_64_T_3[6:0] ? myVec_35 : _GEN_8268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8270 = 7'h24 == _myNewVec_64_T_3[6:0] ? myVec_36 : _GEN_8269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8271 = 7'h25 == _myNewVec_64_T_3[6:0] ? myVec_37 : _GEN_8270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8272 = 7'h26 == _myNewVec_64_T_3[6:0] ? myVec_38 : _GEN_8271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8273 = 7'h27 == _myNewVec_64_T_3[6:0] ? myVec_39 : _GEN_8272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8274 = 7'h28 == _myNewVec_64_T_3[6:0] ? myVec_40 : _GEN_8273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8275 = 7'h29 == _myNewVec_64_T_3[6:0] ? myVec_41 : _GEN_8274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8276 = 7'h2a == _myNewVec_64_T_3[6:0] ? myVec_42 : _GEN_8275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8277 = 7'h2b == _myNewVec_64_T_3[6:0] ? myVec_43 : _GEN_8276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8278 = 7'h2c == _myNewVec_64_T_3[6:0] ? myVec_44 : _GEN_8277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8279 = 7'h2d == _myNewVec_64_T_3[6:0] ? myVec_45 : _GEN_8278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8280 = 7'h2e == _myNewVec_64_T_3[6:0] ? myVec_46 : _GEN_8279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8281 = 7'h2f == _myNewVec_64_T_3[6:0] ? myVec_47 : _GEN_8280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8282 = 7'h30 == _myNewVec_64_T_3[6:0] ? myVec_48 : _GEN_8281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8283 = 7'h31 == _myNewVec_64_T_3[6:0] ? myVec_49 : _GEN_8282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8284 = 7'h32 == _myNewVec_64_T_3[6:0] ? myVec_50 : _GEN_8283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8285 = 7'h33 == _myNewVec_64_T_3[6:0] ? myVec_51 : _GEN_8284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8286 = 7'h34 == _myNewVec_64_T_3[6:0] ? myVec_52 : _GEN_8285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8287 = 7'h35 == _myNewVec_64_T_3[6:0] ? myVec_53 : _GEN_8286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8288 = 7'h36 == _myNewVec_64_T_3[6:0] ? myVec_54 : _GEN_8287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8289 = 7'h37 == _myNewVec_64_T_3[6:0] ? myVec_55 : _GEN_8288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8290 = 7'h38 == _myNewVec_64_T_3[6:0] ? myVec_56 : _GEN_8289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8291 = 7'h39 == _myNewVec_64_T_3[6:0] ? myVec_57 : _GEN_8290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8292 = 7'h3a == _myNewVec_64_T_3[6:0] ? myVec_58 : _GEN_8291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8293 = 7'h3b == _myNewVec_64_T_3[6:0] ? myVec_59 : _GEN_8292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8294 = 7'h3c == _myNewVec_64_T_3[6:0] ? myVec_60 : _GEN_8293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8295 = 7'h3d == _myNewVec_64_T_3[6:0] ? myVec_61 : _GEN_8294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8296 = 7'h3e == _myNewVec_64_T_3[6:0] ? myVec_62 : _GEN_8295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8297 = 7'h3f == _myNewVec_64_T_3[6:0] ? myVec_63 : _GEN_8296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8298 = 7'h40 == _myNewVec_64_T_3[6:0] ? myVec_64 : _GEN_8297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8299 = 7'h41 == _myNewVec_64_T_3[6:0] ? myVec_65 : _GEN_8298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8300 = 7'h42 == _myNewVec_64_T_3[6:0] ? myVec_66 : _GEN_8299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8301 = 7'h43 == _myNewVec_64_T_3[6:0] ? myVec_67 : _GEN_8300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8302 = 7'h44 == _myNewVec_64_T_3[6:0] ? myVec_68 : _GEN_8301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8303 = 7'h45 == _myNewVec_64_T_3[6:0] ? myVec_69 : _GEN_8302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8304 = 7'h46 == _myNewVec_64_T_3[6:0] ? myVec_70 : _GEN_8303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8305 = 7'h47 == _myNewVec_64_T_3[6:0] ? myVec_71 : _GEN_8304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8306 = 7'h48 == _myNewVec_64_T_3[6:0] ? myVec_72 : _GEN_8305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8307 = 7'h49 == _myNewVec_64_T_3[6:0] ? myVec_73 : _GEN_8306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8308 = 7'h4a == _myNewVec_64_T_3[6:0] ? myVec_74 : _GEN_8307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8309 = 7'h4b == _myNewVec_64_T_3[6:0] ? myVec_75 : _GEN_8308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8310 = 7'h4c == _myNewVec_64_T_3[6:0] ? myVec_76 : _GEN_8309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8311 = 7'h4d == _myNewVec_64_T_3[6:0] ? myVec_77 : _GEN_8310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8312 = 7'h4e == _myNewVec_64_T_3[6:0] ? myVec_78 : _GEN_8311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8313 = 7'h4f == _myNewVec_64_T_3[6:0] ? myVec_79 : _GEN_8312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8314 = 7'h50 == _myNewVec_64_T_3[6:0] ? myVec_80 : _GEN_8313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8315 = 7'h51 == _myNewVec_64_T_3[6:0] ? myVec_81 : _GEN_8314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8316 = 7'h52 == _myNewVec_64_T_3[6:0] ? myVec_82 : _GEN_8315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8317 = 7'h53 == _myNewVec_64_T_3[6:0] ? myVec_83 : _GEN_8316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8318 = 7'h54 == _myNewVec_64_T_3[6:0] ? myVec_84 : _GEN_8317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8319 = 7'h55 == _myNewVec_64_T_3[6:0] ? myVec_85 : _GEN_8318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8320 = 7'h56 == _myNewVec_64_T_3[6:0] ? myVec_86 : _GEN_8319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8321 = 7'h57 == _myNewVec_64_T_3[6:0] ? myVec_87 : _GEN_8320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8322 = 7'h58 == _myNewVec_64_T_3[6:0] ? myVec_88 : _GEN_8321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8323 = 7'h59 == _myNewVec_64_T_3[6:0] ? myVec_89 : _GEN_8322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8324 = 7'h5a == _myNewVec_64_T_3[6:0] ? myVec_90 : _GEN_8323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8325 = 7'h5b == _myNewVec_64_T_3[6:0] ? myVec_91 : _GEN_8324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8326 = 7'h5c == _myNewVec_64_T_3[6:0] ? myVec_92 : _GEN_8325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8327 = 7'h5d == _myNewVec_64_T_3[6:0] ? myVec_93 : _GEN_8326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8328 = 7'h5e == _myNewVec_64_T_3[6:0] ? myVec_94 : _GEN_8327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8329 = 7'h5f == _myNewVec_64_T_3[6:0] ? myVec_95 : _GEN_8328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8330 = 7'h60 == _myNewVec_64_T_3[6:0] ? myVec_96 : _GEN_8329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8331 = 7'h61 == _myNewVec_64_T_3[6:0] ? myVec_97 : _GEN_8330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8332 = 7'h62 == _myNewVec_64_T_3[6:0] ? myVec_98 : _GEN_8331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8333 = 7'h63 == _myNewVec_64_T_3[6:0] ? myVec_99 : _GEN_8332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8334 = 7'h64 == _myNewVec_64_T_3[6:0] ? myVec_100 : _GEN_8333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8335 = 7'h65 == _myNewVec_64_T_3[6:0] ? myVec_101 : _GEN_8334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8336 = 7'h66 == _myNewVec_64_T_3[6:0] ? myVec_102 : _GEN_8335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8337 = 7'h67 == _myNewVec_64_T_3[6:0] ? myVec_103 : _GEN_8336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8338 = 7'h68 == _myNewVec_64_T_3[6:0] ? myVec_104 : _GEN_8337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8339 = 7'h69 == _myNewVec_64_T_3[6:0] ? myVec_105 : _GEN_8338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8340 = 7'h6a == _myNewVec_64_T_3[6:0] ? myVec_106 : _GEN_8339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8341 = 7'h6b == _myNewVec_64_T_3[6:0] ? myVec_107 : _GEN_8340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8342 = 7'h6c == _myNewVec_64_T_3[6:0] ? myVec_108 : _GEN_8341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8343 = 7'h6d == _myNewVec_64_T_3[6:0] ? myVec_109 : _GEN_8342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8344 = 7'h6e == _myNewVec_64_T_3[6:0] ? myVec_110 : _GEN_8343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8345 = 7'h6f == _myNewVec_64_T_3[6:0] ? myVec_111 : _GEN_8344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8346 = 7'h70 == _myNewVec_64_T_3[6:0] ? myVec_112 : _GEN_8345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8347 = 7'h71 == _myNewVec_64_T_3[6:0] ? myVec_113 : _GEN_8346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8348 = 7'h72 == _myNewVec_64_T_3[6:0] ? myVec_114 : _GEN_8347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8349 = 7'h73 == _myNewVec_64_T_3[6:0] ? myVec_115 : _GEN_8348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8350 = 7'h74 == _myNewVec_64_T_3[6:0] ? myVec_116 : _GEN_8349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8351 = 7'h75 == _myNewVec_64_T_3[6:0] ? myVec_117 : _GEN_8350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8352 = 7'h76 == _myNewVec_64_T_3[6:0] ? myVec_118 : _GEN_8351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8353 = 7'h77 == _myNewVec_64_T_3[6:0] ? myVec_119 : _GEN_8352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8354 = 7'h78 == _myNewVec_64_T_3[6:0] ? myVec_120 : _GEN_8353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8355 = 7'h79 == _myNewVec_64_T_3[6:0] ? myVec_121 : _GEN_8354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8356 = 7'h7a == _myNewVec_64_T_3[6:0] ? myVec_122 : _GEN_8355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8357 = 7'h7b == _myNewVec_64_T_3[6:0] ? myVec_123 : _GEN_8356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8358 = 7'h7c == _myNewVec_64_T_3[6:0] ? myVec_124 : _GEN_8357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8359 = 7'h7d == _myNewVec_64_T_3[6:0] ? myVec_125 : _GEN_8358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8360 = 7'h7e == _myNewVec_64_T_3[6:0] ? myVec_126 : _GEN_8359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_64 = 7'h7f == _myNewVec_64_T_3[6:0] ? myVec_127 : _GEN_8360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [255:0] myNewWire_hi_lo_lo_lo = {myNewVec_71,myNewVec_70,myNewVec_69,myNewVec_68,myNewVec_67,myNewVec_66,
    myNewVec_65,myNewVec_64}; // @[hh_datapath_chisel.scala 238:27]
  wire [511:0] myNewWire_hi_lo_lo = {myNewVec_79,myNewVec_78,myNewVec_77,myNewVec_76,myNewVec_75,myNewVec_74,myNewVec_73
    ,myNewVec_72,myNewWire_hi_lo_lo_lo}; // @[hh_datapath_chisel.scala 238:27]
  wire [1023:0] myNewWire_hi_lo = {myNewVec_95,myNewVec_94,myNewVec_93,myNewVec_92,myNewVec_91,myNewVec_90,myNewVec_89,
    myNewVec_88,myNewWire_hi_lo_hi_lo,myNewWire_hi_lo_lo}; // @[hh_datapath_chisel.scala 238:27]
  wire [15:0] _myNewVec_63_T_3 = _myNewVec_127_T_1 + 16'h40; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_8363 = 7'h1 == _myNewVec_63_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8364 = 7'h2 == _myNewVec_63_T_3[6:0] ? myVec_2 : _GEN_8363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8365 = 7'h3 == _myNewVec_63_T_3[6:0] ? myVec_3 : _GEN_8364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8366 = 7'h4 == _myNewVec_63_T_3[6:0] ? myVec_4 : _GEN_8365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8367 = 7'h5 == _myNewVec_63_T_3[6:0] ? myVec_5 : _GEN_8366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8368 = 7'h6 == _myNewVec_63_T_3[6:0] ? myVec_6 : _GEN_8367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8369 = 7'h7 == _myNewVec_63_T_3[6:0] ? myVec_7 : _GEN_8368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8370 = 7'h8 == _myNewVec_63_T_3[6:0] ? myVec_8 : _GEN_8369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8371 = 7'h9 == _myNewVec_63_T_3[6:0] ? myVec_9 : _GEN_8370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8372 = 7'ha == _myNewVec_63_T_3[6:0] ? myVec_10 : _GEN_8371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8373 = 7'hb == _myNewVec_63_T_3[6:0] ? myVec_11 : _GEN_8372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8374 = 7'hc == _myNewVec_63_T_3[6:0] ? myVec_12 : _GEN_8373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8375 = 7'hd == _myNewVec_63_T_3[6:0] ? myVec_13 : _GEN_8374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8376 = 7'he == _myNewVec_63_T_3[6:0] ? myVec_14 : _GEN_8375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8377 = 7'hf == _myNewVec_63_T_3[6:0] ? myVec_15 : _GEN_8376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8378 = 7'h10 == _myNewVec_63_T_3[6:0] ? myVec_16 : _GEN_8377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8379 = 7'h11 == _myNewVec_63_T_3[6:0] ? myVec_17 : _GEN_8378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8380 = 7'h12 == _myNewVec_63_T_3[6:0] ? myVec_18 : _GEN_8379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8381 = 7'h13 == _myNewVec_63_T_3[6:0] ? myVec_19 : _GEN_8380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8382 = 7'h14 == _myNewVec_63_T_3[6:0] ? myVec_20 : _GEN_8381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8383 = 7'h15 == _myNewVec_63_T_3[6:0] ? myVec_21 : _GEN_8382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8384 = 7'h16 == _myNewVec_63_T_3[6:0] ? myVec_22 : _GEN_8383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8385 = 7'h17 == _myNewVec_63_T_3[6:0] ? myVec_23 : _GEN_8384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8386 = 7'h18 == _myNewVec_63_T_3[6:0] ? myVec_24 : _GEN_8385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8387 = 7'h19 == _myNewVec_63_T_3[6:0] ? myVec_25 : _GEN_8386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8388 = 7'h1a == _myNewVec_63_T_3[6:0] ? myVec_26 : _GEN_8387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8389 = 7'h1b == _myNewVec_63_T_3[6:0] ? myVec_27 : _GEN_8388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8390 = 7'h1c == _myNewVec_63_T_3[6:0] ? myVec_28 : _GEN_8389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8391 = 7'h1d == _myNewVec_63_T_3[6:0] ? myVec_29 : _GEN_8390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8392 = 7'h1e == _myNewVec_63_T_3[6:0] ? myVec_30 : _GEN_8391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8393 = 7'h1f == _myNewVec_63_T_3[6:0] ? myVec_31 : _GEN_8392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8394 = 7'h20 == _myNewVec_63_T_3[6:0] ? myVec_32 : _GEN_8393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8395 = 7'h21 == _myNewVec_63_T_3[6:0] ? myVec_33 : _GEN_8394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8396 = 7'h22 == _myNewVec_63_T_3[6:0] ? myVec_34 : _GEN_8395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8397 = 7'h23 == _myNewVec_63_T_3[6:0] ? myVec_35 : _GEN_8396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8398 = 7'h24 == _myNewVec_63_T_3[6:0] ? myVec_36 : _GEN_8397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8399 = 7'h25 == _myNewVec_63_T_3[6:0] ? myVec_37 : _GEN_8398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8400 = 7'h26 == _myNewVec_63_T_3[6:0] ? myVec_38 : _GEN_8399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8401 = 7'h27 == _myNewVec_63_T_3[6:0] ? myVec_39 : _GEN_8400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8402 = 7'h28 == _myNewVec_63_T_3[6:0] ? myVec_40 : _GEN_8401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8403 = 7'h29 == _myNewVec_63_T_3[6:0] ? myVec_41 : _GEN_8402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8404 = 7'h2a == _myNewVec_63_T_3[6:0] ? myVec_42 : _GEN_8403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8405 = 7'h2b == _myNewVec_63_T_3[6:0] ? myVec_43 : _GEN_8404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8406 = 7'h2c == _myNewVec_63_T_3[6:0] ? myVec_44 : _GEN_8405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8407 = 7'h2d == _myNewVec_63_T_3[6:0] ? myVec_45 : _GEN_8406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8408 = 7'h2e == _myNewVec_63_T_3[6:0] ? myVec_46 : _GEN_8407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8409 = 7'h2f == _myNewVec_63_T_3[6:0] ? myVec_47 : _GEN_8408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8410 = 7'h30 == _myNewVec_63_T_3[6:0] ? myVec_48 : _GEN_8409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8411 = 7'h31 == _myNewVec_63_T_3[6:0] ? myVec_49 : _GEN_8410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8412 = 7'h32 == _myNewVec_63_T_3[6:0] ? myVec_50 : _GEN_8411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8413 = 7'h33 == _myNewVec_63_T_3[6:0] ? myVec_51 : _GEN_8412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8414 = 7'h34 == _myNewVec_63_T_3[6:0] ? myVec_52 : _GEN_8413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8415 = 7'h35 == _myNewVec_63_T_3[6:0] ? myVec_53 : _GEN_8414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8416 = 7'h36 == _myNewVec_63_T_3[6:0] ? myVec_54 : _GEN_8415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8417 = 7'h37 == _myNewVec_63_T_3[6:0] ? myVec_55 : _GEN_8416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8418 = 7'h38 == _myNewVec_63_T_3[6:0] ? myVec_56 : _GEN_8417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8419 = 7'h39 == _myNewVec_63_T_3[6:0] ? myVec_57 : _GEN_8418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8420 = 7'h3a == _myNewVec_63_T_3[6:0] ? myVec_58 : _GEN_8419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8421 = 7'h3b == _myNewVec_63_T_3[6:0] ? myVec_59 : _GEN_8420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8422 = 7'h3c == _myNewVec_63_T_3[6:0] ? myVec_60 : _GEN_8421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8423 = 7'h3d == _myNewVec_63_T_3[6:0] ? myVec_61 : _GEN_8422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8424 = 7'h3e == _myNewVec_63_T_3[6:0] ? myVec_62 : _GEN_8423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8425 = 7'h3f == _myNewVec_63_T_3[6:0] ? myVec_63 : _GEN_8424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8426 = 7'h40 == _myNewVec_63_T_3[6:0] ? myVec_64 : _GEN_8425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8427 = 7'h41 == _myNewVec_63_T_3[6:0] ? myVec_65 : _GEN_8426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8428 = 7'h42 == _myNewVec_63_T_3[6:0] ? myVec_66 : _GEN_8427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8429 = 7'h43 == _myNewVec_63_T_3[6:0] ? myVec_67 : _GEN_8428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8430 = 7'h44 == _myNewVec_63_T_3[6:0] ? myVec_68 : _GEN_8429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8431 = 7'h45 == _myNewVec_63_T_3[6:0] ? myVec_69 : _GEN_8430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8432 = 7'h46 == _myNewVec_63_T_3[6:0] ? myVec_70 : _GEN_8431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8433 = 7'h47 == _myNewVec_63_T_3[6:0] ? myVec_71 : _GEN_8432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8434 = 7'h48 == _myNewVec_63_T_3[6:0] ? myVec_72 : _GEN_8433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8435 = 7'h49 == _myNewVec_63_T_3[6:0] ? myVec_73 : _GEN_8434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8436 = 7'h4a == _myNewVec_63_T_3[6:0] ? myVec_74 : _GEN_8435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8437 = 7'h4b == _myNewVec_63_T_3[6:0] ? myVec_75 : _GEN_8436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8438 = 7'h4c == _myNewVec_63_T_3[6:0] ? myVec_76 : _GEN_8437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8439 = 7'h4d == _myNewVec_63_T_3[6:0] ? myVec_77 : _GEN_8438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8440 = 7'h4e == _myNewVec_63_T_3[6:0] ? myVec_78 : _GEN_8439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8441 = 7'h4f == _myNewVec_63_T_3[6:0] ? myVec_79 : _GEN_8440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8442 = 7'h50 == _myNewVec_63_T_3[6:0] ? myVec_80 : _GEN_8441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8443 = 7'h51 == _myNewVec_63_T_3[6:0] ? myVec_81 : _GEN_8442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8444 = 7'h52 == _myNewVec_63_T_3[6:0] ? myVec_82 : _GEN_8443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8445 = 7'h53 == _myNewVec_63_T_3[6:0] ? myVec_83 : _GEN_8444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8446 = 7'h54 == _myNewVec_63_T_3[6:0] ? myVec_84 : _GEN_8445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8447 = 7'h55 == _myNewVec_63_T_3[6:0] ? myVec_85 : _GEN_8446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8448 = 7'h56 == _myNewVec_63_T_3[6:0] ? myVec_86 : _GEN_8447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8449 = 7'h57 == _myNewVec_63_T_3[6:0] ? myVec_87 : _GEN_8448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8450 = 7'h58 == _myNewVec_63_T_3[6:0] ? myVec_88 : _GEN_8449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8451 = 7'h59 == _myNewVec_63_T_3[6:0] ? myVec_89 : _GEN_8450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8452 = 7'h5a == _myNewVec_63_T_3[6:0] ? myVec_90 : _GEN_8451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8453 = 7'h5b == _myNewVec_63_T_3[6:0] ? myVec_91 : _GEN_8452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8454 = 7'h5c == _myNewVec_63_T_3[6:0] ? myVec_92 : _GEN_8453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8455 = 7'h5d == _myNewVec_63_T_3[6:0] ? myVec_93 : _GEN_8454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8456 = 7'h5e == _myNewVec_63_T_3[6:0] ? myVec_94 : _GEN_8455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8457 = 7'h5f == _myNewVec_63_T_3[6:0] ? myVec_95 : _GEN_8456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8458 = 7'h60 == _myNewVec_63_T_3[6:0] ? myVec_96 : _GEN_8457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8459 = 7'h61 == _myNewVec_63_T_3[6:0] ? myVec_97 : _GEN_8458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8460 = 7'h62 == _myNewVec_63_T_3[6:0] ? myVec_98 : _GEN_8459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8461 = 7'h63 == _myNewVec_63_T_3[6:0] ? myVec_99 : _GEN_8460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8462 = 7'h64 == _myNewVec_63_T_3[6:0] ? myVec_100 : _GEN_8461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8463 = 7'h65 == _myNewVec_63_T_3[6:0] ? myVec_101 : _GEN_8462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8464 = 7'h66 == _myNewVec_63_T_3[6:0] ? myVec_102 : _GEN_8463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8465 = 7'h67 == _myNewVec_63_T_3[6:0] ? myVec_103 : _GEN_8464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8466 = 7'h68 == _myNewVec_63_T_3[6:0] ? myVec_104 : _GEN_8465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8467 = 7'h69 == _myNewVec_63_T_3[6:0] ? myVec_105 : _GEN_8466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8468 = 7'h6a == _myNewVec_63_T_3[6:0] ? myVec_106 : _GEN_8467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8469 = 7'h6b == _myNewVec_63_T_3[6:0] ? myVec_107 : _GEN_8468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8470 = 7'h6c == _myNewVec_63_T_3[6:0] ? myVec_108 : _GEN_8469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8471 = 7'h6d == _myNewVec_63_T_3[6:0] ? myVec_109 : _GEN_8470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8472 = 7'h6e == _myNewVec_63_T_3[6:0] ? myVec_110 : _GEN_8471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8473 = 7'h6f == _myNewVec_63_T_3[6:0] ? myVec_111 : _GEN_8472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8474 = 7'h70 == _myNewVec_63_T_3[6:0] ? myVec_112 : _GEN_8473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8475 = 7'h71 == _myNewVec_63_T_3[6:0] ? myVec_113 : _GEN_8474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8476 = 7'h72 == _myNewVec_63_T_3[6:0] ? myVec_114 : _GEN_8475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8477 = 7'h73 == _myNewVec_63_T_3[6:0] ? myVec_115 : _GEN_8476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8478 = 7'h74 == _myNewVec_63_T_3[6:0] ? myVec_116 : _GEN_8477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8479 = 7'h75 == _myNewVec_63_T_3[6:0] ? myVec_117 : _GEN_8478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8480 = 7'h76 == _myNewVec_63_T_3[6:0] ? myVec_118 : _GEN_8479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8481 = 7'h77 == _myNewVec_63_T_3[6:0] ? myVec_119 : _GEN_8480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8482 = 7'h78 == _myNewVec_63_T_3[6:0] ? myVec_120 : _GEN_8481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8483 = 7'h79 == _myNewVec_63_T_3[6:0] ? myVec_121 : _GEN_8482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8484 = 7'h7a == _myNewVec_63_T_3[6:0] ? myVec_122 : _GEN_8483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8485 = 7'h7b == _myNewVec_63_T_3[6:0] ? myVec_123 : _GEN_8484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8486 = 7'h7c == _myNewVec_63_T_3[6:0] ? myVec_124 : _GEN_8485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8487 = 7'h7d == _myNewVec_63_T_3[6:0] ? myVec_125 : _GEN_8486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8488 = 7'h7e == _myNewVec_63_T_3[6:0] ? myVec_126 : _GEN_8487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_63 = 7'h7f == _myNewVec_63_T_3[6:0] ? myVec_127 : _GEN_8488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_62_T_3 = _myNewVec_127_T_1 + 16'h41; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_8491 = 7'h1 == _myNewVec_62_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8492 = 7'h2 == _myNewVec_62_T_3[6:0] ? myVec_2 : _GEN_8491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8493 = 7'h3 == _myNewVec_62_T_3[6:0] ? myVec_3 : _GEN_8492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8494 = 7'h4 == _myNewVec_62_T_3[6:0] ? myVec_4 : _GEN_8493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8495 = 7'h5 == _myNewVec_62_T_3[6:0] ? myVec_5 : _GEN_8494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8496 = 7'h6 == _myNewVec_62_T_3[6:0] ? myVec_6 : _GEN_8495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8497 = 7'h7 == _myNewVec_62_T_3[6:0] ? myVec_7 : _GEN_8496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8498 = 7'h8 == _myNewVec_62_T_3[6:0] ? myVec_8 : _GEN_8497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8499 = 7'h9 == _myNewVec_62_T_3[6:0] ? myVec_9 : _GEN_8498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8500 = 7'ha == _myNewVec_62_T_3[6:0] ? myVec_10 : _GEN_8499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8501 = 7'hb == _myNewVec_62_T_3[6:0] ? myVec_11 : _GEN_8500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8502 = 7'hc == _myNewVec_62_T_3[6:0] ? myVec_12 : _GEN_8501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8503 = 7'hd == _myNewVec_62_T_3[6:0] ? myVec_13 : _GEN_8502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8504 = 7'he == _myNewVec_62_T_3[6:0] ? myVec_14 : _GEN_8503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8505 = 7'hf == _myNewVec_62_T_3[6:0] ? myVec_15 : _GEN_8504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8506 = 7'h10 == _myNewVec_62_T_3[6:0] ? myVec_16 : _GEN_8505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8507 = 7'h11 == _myNewVec_62_T_3[6:0] ? myVec_17 : _GEN_8506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8508 = 7'h12 == _myNewVec_62_T_3[6:0] ? myVec_18 : _GEN_8507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8509 = 7'h13 == _myNewVec_62_T_3[6:0] ? myVec_19 : _GEN_8508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8510 = 7'h14 == _myNewVec_62_T_3[6:0] ? myVec_20 : _GEN_8509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8511 = 7'h15 == _myNewVec_62_T_3[6:0] ? myVec_21 : _GEN_8510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8512 = 7'h16 == _myNewVec_62_T_3[6:0] ? myVec_22 : _GEN_8511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8513 = 7'h17 == _myNewVec_62_T_3[6:0] ? myVec_23 : _GEN_8512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8514 = 7'h18 == _myNewVec_62_T_3[6:0] ? myVec_24 : _GEN_8513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8515 = 7'h19 == _myNewVec_62_T_3[6:0] ? myVec_25 : _GEN_8514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8516 = 7'h1a == _myNewVec_62_T_3[6:0] ? myVec_26 : _GEN_8515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8517 = 7'h1b == _myNewVec_62_T_3[6:0] ? myVec_27 : _GEN_8516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8518 = 7'h1c == _myNewVec_62_T_3[6:0] ? myVec_28 : _GEN_8517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8519 = 7'h1d == _myNewVec_62_T_3[6:0] ? myVec_29 : _GEN_8518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8520 = 7'h1e == _myNewVec_62_T_3[6:0] ? myVec_30 : _GEN_8519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8521 = 7'h1f == _myNewVec_62_T_3[6:0] ? myVec_31 : _GEN_8520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8522 = 7'h20 == _myNewVec_62_T_3[6:0] ? myVec_32 : _GEN_8521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8523 = 7'h21 == _myNewVec_62_T_3[6:0] ? myVec_33 : _GEN_8522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8524 = 7'h22 == _myNewVec_62_T_3[6:0] ? myVec_34 : _GEN_8523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8525 = 7'h23 == _myNewVec_62_T_3[6:0] ? myVec_35 : _GEN_8524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8526 = 7'h24 == _myNewVec_62_T_3[6:0] ? myVec_36 : _GEN_8525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8527 = 7'h25 == _myNewVec_62_T_3[6:0] ? myVec_37 : _GEN_8526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8528 = 7'h26 == _myNewVec_62_T_3[6:0] ? myVec_38 : _GEN_8527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8529 = 7'h27 == _myNewVec_62_T_3[6:0] ? myVec_39 : _GEN_8528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8530 = 7'h28 == _myNewVec_62_T_3[6:0] ? myVec_40 : _GEN_8529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8531 = 7'h29 == _myNewVec_62_T_3[6:0] ? myVec_41 : _GEN_8530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8532 = 7'h2a == _myNewVec_62_T_3[6:0] ? myVec_42 : _GEN_8531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8533 = 7'h2b == _myNewVec_62_T_3[6:0] ? myVec_43 : _GEN_8532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8534 = 7'h2c == _myNewVec_62_T_3[6:0] ? myVec_44 : _GEN_8533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8535 = 7'h2d == _myNewVec_62_T_3[6:0] ? myVec_45 : _GEN_8534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8536 = 7'h2e == _myNewVec_62_T_3[6:0] ? myVec_46 : _GEN_8535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8537 = 7'h2f == _myNewVec_62_T_3[6:0] ? myVec_47 : _GEN_8536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8538 = 7'h30 == _myNewVec_62_T_3[6:0] ? myVec_48 : _GEN_8537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8539 = 7'h31 == _myNewVec_62_T_3[6:0] ? myVec_49 : _GEN_8538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8540 = 7'h32 == _myNewVec_62_T_3[6:0] ? myVec_50 : _GEN_8539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8541 = 7'h33 == _myNewVec_62_T_3[6:0] ? myVec_51 : _GEN_8540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8542 = 7'h34 == _myNewVec_62_T_3[6:0] ? myVec_52 : _GEN_8541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8543 = 7'h35 == _myNewVec_62_T_3[6:0] ? myVec_53 : _GEN_8542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8544 = 7'h36 == _myNewVec_62_T_3[6:0] ? myVec_54 : _GEN_8543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8545 = 7'h37 == _myNewVec_62_T_3[6:0] ? myVec_55 : _GEN_8544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8546 = 7'h38 == _myNewVec_62_T_3[6:0] ? myVec_56 : _GEN_8545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8547 = 7'h39 == _myNewVec_62_T_3[6:0] ? myVec_57 : _GEN_8546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8548 = 7'h3a == _myNewVec_62_T_3[6:0] ? myVec_58 : _GEN_8547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8549 = 7'h3b == _myNewVec_62_T_3[6:0] ? myVec_59 : _GEN_8548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8550 = 7'h3c == _myNewVec_62_T_3[6:0] ? myVec_60 : _GEN_8549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8551 = 7'h3d == _myNewVec_62_T_3[6:0] ? myVec_61 : _GEN_8550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8552 = 7'h3e == _myNewVec_62_T_3[6:0] ? myVec_62 : _GEN_8551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8553 = 7'h3f == _myNewVec_62_T_3[6:0] ? myVec_63 : _GEN_8552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8554 = 7'h40 == _myNewVec_62_T_3[6:0] ? myVec_64 : _GEN_8553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8555 = 7'h41 == _myNewVec_62_T_3[6:0] ? myVec_65 : _GEN_8554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8556 = 7'h42 == _myNewVec_62_T_3[6:0] ? myVec_66 : _GEN_8555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8557 = 7'h43 == _myNewVec_62_T_3[6:0] ? myVec_67 : _GEN_8556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8558 = 7'h44 == _myNewVec_62_T_3[6:0] ? myVec_68 : _GEN_8557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8559 = 7'h45 == _myNewVec_62_T_3[6:0] ? myVec_69 : _GEN_8558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8560 = 7'h46 == _myNewVec_62_T_3[6:0] ? myVec_70 : _GEN_8559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8561 = 7'h47 == _myNewVec_62_T_3[6:0] ? myVec_71 : _GEN_8560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8562 = 7'h48 == _myNewVec_62_T_3[6:0] ? myVec_72 : _GEN_8561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8563 = 7'h49 == _myNewVec_62_T_3[6:0] ? myVec_73 : _GEN_8562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8564 = 7'h4a == _myNewVec_62_T_3[6:0] ? myVec_74 : _GEN_8563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8565 = 7'h4b == _myNewVec_62_T_3[6:0] ? myVec_75 : _GEN_8564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8566 = 7'h4c == _myNewVec_62_T_3[6:0] ? myVec_76 : _GEN_8565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8567 = 7'h4d == _myNewVec_62_T_3[6:0] ? myVec_77 : _GEN_8566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8568 = 7'h4e == _myNewVec_62_T_3[6:0] ? myVec_78 : _GEN_8567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8569 = 7'h4f == _myNewVec_62_T_3[6:0] ? myVec_79 : _GEN_8568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8570 = 7'h50 == _myNewVec_62_T_3[6:0] ? myVec_80 : _GEN_8569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8571 = 7'h51 == _myNewVec_62_T_3[6:0] ? myVec_81 : _GEN_8570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8572 = 7'h52 == _myNewVec_62_T_3[6:0] ? myVec_82 : _GEN_8571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8573 = 7'h53 == _myNewVec_62_T_3[6:0] ? myVec_83 : _GEN_8572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8574 = 7'h54 == _myNewVec_62_T_3[6:0] ? myVec_84 : _GEN_8573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8575 = 7'h55 == _myNewVec_62_T_3[6:0] ? myVec_85 : _GEN_8574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8576 = 7'h56 == _myNewVec_62_T_3[6:0] ? myVec_86 : _GEN_8575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8577 = 7'h57 == _myNewVec_62_T_3[6:0] ? myVec_87 : _GEN_8576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8578 = 7'h58 == _myNewVec_62_T_3[6:0] ? myVec_88 : _GEN_8577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8579 = 7'h59 == _myNewVec_62_T_3[6:0] ? myVec_89 : _GEN_8578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8580 = 7'h5a == _myNewVec_62_T_3[6:0] ? myVec_90 : _GEN_8579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8581 = 7'h5b == _myNewVec_62_T_3[6:0] ? myVec_91 : _GEN_8580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8582 = 7'h5c == _myNewVec_62_T_3[6:0] ? myVec_92 : _GEN_8581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8583 = 7'h5d == _myNewVec_62_T_3[6:0] ? myVec_93 : _GEN_8582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8584 = 7'h5e == _myNewVec_62_T_3[6:0] ? myVec_94 : _GEN_8583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8585 = 7'h5f == _myNewVec_62_T_3[6:0] ? myVec_95 : _GEN_8584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8586 = 7'h60 == _myNewVec_62_T_3[6:0] ? myVec_96 : _GEN_8585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8587 = 7'h61 == _myNewVec_62_T_3[6:0] ? myVec_97 : _GEN_8586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8588 = 7'h62 == _myNewVec_62_T_3[6:0] ? myVec_98 : _GEN_8587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8589 = 7'h63 == _myNewVec_62_T_3[6:0] ? myVec_99 : _GEN_8588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8590 = 7'h64 == _myNewVec_62_T_3[6:0] ? myVec_100 : _GEN_8589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8591 = 7'h65 == _myNewVec_62_T_3[6:0] ? myVec_101 : _GEN_8590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8592 = 7'h66 == _myNewVec_62_T_3[6:0] ? myVec_102 : _GEN_8591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8593 = 7'h67 == _myNewVec_62_T_3[6:0] ? myVec_103 : _GEN_8592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8594 = 7'h68 == _myNewVec_62_T_3[6:0] ? myVec_104 : _GEN_8593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8595 = 7'h69 == _myNewVec_62_T_3[6:0] ? myVec_105 : _GEN_8594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8596 = 7'h6a == _myNewVec_62_T_3[6:0] ? myVec_106 : _GEN_8595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8597 = 7'h6b == _myNewVec_62_T_3[6:0] ? myVec_107 : _GEN_8596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8598 = 7'h6c == _myNewVec_62_T_3[6:0] ? myVec_108 : _GEN_8597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8599 = 7'h6d == _myNewVec_62_T_3[6:0] ? myVec_109 : _GEN_8598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8600 = 7'h6e == _myNewVec_62_T_3[6:0] ? myVec_110 : _GEN_8599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8601 = 7'h6f == _myNewVec_62_T_3[6:0] ? myVec_111 : _GEN_8600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8602 = 7'h70 == _myNewVec_62_T_3[6:0] ? myVec_112 : _GEN_8601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8603 = 7'h71 == _myNewVec_62_T_3[6:0] ? myVec_113 : _GEN_8602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8604 = 7'h72 == _myNewVec_62_T_3[6:0] ? myVec_114 : _GEN_8603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8605 = 7'h73 == _myNewVec_62_T_3[6:0] ? myVec_115 : _GEN_8604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8606 = 7'h74 == _myNewVec_62_T_3[6:0] ? myVec_116 : _GEN_8605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8607 = 7'h75 == _myNewVec_62_T_3[6:0] ? myVec_117 : _GEN_8606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8608 = 7'h76 == _myNewVec_62_T_3[6:0] ? myVec_118 : _GEN_8607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8609 = 7'h77 == _myNewVec_62_T_3[6:0] ? myVec_119 : _GEN_8608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8610 = 7'h78 == _myNewVec_62_T_3[6:0] ? myVec_120 : _GEN_8609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8611 = 7'h79 == _myNewVec_62_T_3[6:0] ? myVec_121 : _GEN_8610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8612 = 7'h7a == _myNewVec_62_T_3[6:0] ? myVec_122 : _GEN_8611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8613 = 7'h7b == _myNewVec_62_T_3[6:0] ? myVec_123 : _GEN_8612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8614 = 7'h7c == _myNewVec_62_T_3[6:0] ? myVec_124 : _GEN_8613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8615 = 7'h7d == _myNewVec_62_T_3[6:0] ? myVec_125 : _GEN_8614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8616 = 7'h7e == _myNewVec_62_T_3[6:0] ? myVec_126 : _GEN_8615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_62 = 7'h7f == _myNewVec_62_T_3[6:0] ? myVec_127 : _GEN_8616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_61_T_3 = _myNewVec_127_T_1 + 16'h42; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_8619 = 7'h1 == _myNewVec_61_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8620 = 7'h2 == _myNewVec_61_T_3[6:0] ? myVec_2 : _GEN_8619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8621 = 7'h3 == _myNewVec_61_T_3[6:0] ? myVec_3 : _GEN_8620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8622 = 7'h4 == _myNewVec_61_T_3[6:0] ? myVec_4 : _GEN_8621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8623 = 7'h5 == _myNewVec_61_T_3[6:0] ? myVec_5 : _GEN_8622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8624 = 7'h6 == _myNewVec_61_T_3[6:0] ? myVec_6 : _GEN_8623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8625 = 7'h7 == _myNewVec_61_T_3[6:0] ? myVec_7 : _GEN_8624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8626 = 7'h8 == _myNewVec_61_T_3[6:0] ? myVec_8 : _GEN_8625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8627 = 7'h9 == _myNewVec_61_T_3[6:0] ? myVec_9 : _GEN_8626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8628 = 7'ha == _myNewVec_61_T_3[6:0] ? myVec_10 : _GEN_8627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8629 = 7'hb == _myNewVec_61_T_3[6:0] ? myVec_11 : _GEN_8628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8630 = 7'hc == _myNewVec_61_T_3[6:0] ? myVec_12 : _GEN_8629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8631 = 7'hd == _myNewVec_61_T_3[6:0] ? myVec_13 : _GEN_8630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8632 = 7'he == _myNewVec_61_T_3[6:0] ? myVec_14 : _GEN_8631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8633 = 7'hf == _myNewVec_61_T_3[6:0] ? myVec_15 : _GEN_8632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8634 = 7'h10 == _myNewVec_61_T_3[6:0] ? myVec_16 : _GEN_8633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8635 = 7'h11 == _myNewVec_61_T_3[6:0] ? myVec_17 : _GEN_8634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8636 = 7'h12 == _myNewVec_61_T_3[6:0] ? myVec_18 : _GEN_8635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8637 = 7'h13 == _myNewVec_61_T_3[6:0] ? myVec_19 : _GEN_8636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8638 = 7'h14 == _myNewVec_61_T_3[6:0] ? myVec_20 : _GEN_8637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8639 = 7'h15 == _myNewVec_61_T_3[6:0] ? myVec_21 : _GEN_8638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8640 = 7'h16 == _myNewVec_61_T_3[6:0] ? myVec_22 : _GEN_8639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8641 = 7'h17 == _myNewVec_61_T_3[6:0] ? myVec_23 : _GEN_8640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8642 = 7'h18 == _myNewVec_61_T_3[6:0] ? myVec_24 : _GEN_8641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8643 = 7'h19 == _myNewVec_61_T_3[6:0] ? myVec_25 : _GEN_8642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8644 = 7'h1a == _myNewVec_61_T_3[6:0] ? myVec_26 : _GEN_8643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8645 = 7'h1b == _myNewVec_61_T_3[6:0] ? myVec_27 : _GEN_8644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8646 = 7'h1c == _myNewVec_61_T_3[6:0] ? myVec_28 : _GEN_8645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8647 = 7'h1d == _myNewVec_61_T_3[6:0] ? myVec_29 : _GEN_8646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8648 = 7'h1e == _myNewVec_61_T_3[6:0] ? myVec_30 : _GEN_8647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8649 = 7'h1f == _myNewVec_61_T_3[6:0] ? myVec_31 : _GEN_8648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8650 = 7'h20 == _myNewVec_61_T_3[6:0] ? myVec_32 : _GEN_8649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8651 = 7'h21 == _myNewVec_61_T_3[6:0] ? myVec_33 : _GEN_8650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8652 = 7'h22 == _myNewVec_61_T_3[6:0] ? myVec_34 : _GEN_8651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8653 = 7'h23 == _myNewVec_61_T_3[6:0] ? myVec_35 : _GEN_8652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8654 = 7'h24 == _myNewVec_61_T_3[6:0] ? myVec_36 : _GEN_8653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8655 = 7'h25 == _myNewVec_61_T_3[6:0] ? myVec_37 : _GEN_8654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8656 = 7'h26 == _myNewVec_61_T_3[6:0] ? myVec_38 : _GEN_8655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8657 = 7'h27 == _myNewVec_61_T_3[6:0] ? myVec_39 : _GEN_8656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8658 = 7'h28 == _myNewVec_61_T_3[6:0] ? myVec_40 : _GEN_8657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8659 = 7'h29 == _myNewVec_61_T_3[6:0] ? myVec_41 : _GEN_8658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8660 = 7'h2a == _myNewVec_61_T_3[6:0] ? myVec_42 : _GEN_8659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8661 = 7'h2b == _myNewVec_61_T_3[6:0] ? myVec_43 : _GEN_8660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8662 = 7'h2c == _myNewVec_61_T_3[6:0] ? myVec_44 : _GEN_8661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8663 = 7'h2d == _myNewVec_61_T_3[6:0] ? myVec_45 : _GEN_8662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8664 = 7'h2e == _myNewVec_61_T_3[6:0] ? myVec_46 : _GEN_8663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8665 = 7'h2f == _myNewVec_61_T_3[6:0] ? myVec_47 : _GEN_8664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8666 = 7'h30 == _myNewVec_61_T_3[6:0] ? myVec_48 : _GEN_8665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8667 = 7'h31 == _myNewVec_61_T_3[6:0] ? myVec_49 : _GEN_8666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8668 = 7'h32 == _myNewVec_61_T_3[6:0] ? myVec_50 : _GEN_8667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8669 = 7'h33 == _myNewVec_61_T_3[6:0] ? myVec_51 : _GEN_8668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8670 = 7'h34 == _myNewVec_61_T_3[6:0] ? myVec_52 : _GEN_8669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8671 = 7'h35 == _myNewVec_61_T_3[6:0] ? myVec_53 : _GEN_8670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8672 = 7'h36 == _myNewVec_61_T_3[6:0] ? myVec_54 : _GEN_8671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8673 = 7'h37 == _myNewVec_61_T_3[6:0] ? myVec_55 : _GEN_8672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8674 = 7'h38 == _myNewVec_61_T_3[6:0] ? myVec_56 : _GEN_8673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8675 = 7'h39 == _myNewVec_61_T_3[6:0] ? myVec_57 : _GEN_8674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8676 = 7'h3a == _myNewVec_61_T_3[6:0] ? myVec_58 : _GEN_8675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8677 = 7'h3b == _myNewVec_61_T_3[6:0] ? myVec_59 : _GEN_8676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8678 = 7'h3c == _myNewVec_61_T_3[6:0] ? myVec_60 : _GEN_8677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8679 = 7'h3d == _myNewVec_61_T_3[6:0] ? myVec_61 : _GEN_8678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8680 = 7'h3e == _myNewVec_61_T_3[6:0] ? myVec_62 : _GEN_8679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8681 = 7'h3f == _myNewVec_61_T_3[6:0] ? myVec_63 : _GEN_8680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8682 = 7'h40 == _myNewVec_61_T_3[6:0] ? myVec_64 : _GEN_8681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8683 = 7'h41 == _myNewVec_61_T_3[6:0] ? myVec_65 : _GEN_8682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8684 = 7'h42 == _myNewVec_61_T_3[6:0] ? myVec_66 : _GEN_8683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8685 = 7'h43 == _myNewVec_61_T_3[6:0] ? myVec_67 : _GEN_8684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8686 = 7'h44 == _myNewVec_61_T_3[6:0] ? myVec_68 : _GEN_8685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8687 = 7'h45 == _myNewVec_61_T_3[6:0] ? myVec_69 : _GEN_8686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8688 = 7'h46 == _myNewVec_61_T_3[6:0] ? myVec_70 : _GEN_8687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8689 = 7'h47 == _myNewVec_61_T_3[6:0] ? myVec_71 : _GEN_8688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8690 = 7'h48 == _myNewVec_61_T_3[6:0] ? myVec_72 : _GEN_8689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8691 = 7'h49 == _myNewVec_61_T_3[6:0] ? myVec_73 : _GEN_8690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8692 = 7'h4a == _myNewVec_61_T_3[6:0] ? myVec_74 : _GEN_8691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8693 = 7'h4b == _myNewVec_61_T_3[6:0] ? myVec_75 : _GEN_8692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8694 = 7'h4c == _myNewVec_61_T_3[6:0] ? myVec_76 : _GEN_8693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8695 = 7'h4d == _myNewVec_61_T_3[6:0] ? myVec_77 : _GEN_8694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8696 = 7'h4e == _myNewVec_61_T_3[6:0] ? myVec_78 : _GEN_8695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8697 = 7'h4f == _myNewVec_61_T_3[6:0] ? myVec_79 : _GEN_8696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8698 = 7'h50 == _myNewVec_61_T_3[6:0] ? myVec_80 : _GEN_8697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8699 = 7'h51 == _myNewVec_61_T_3[6:0] ? myVec_81 : _GEN_8698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8700 = 7'h52 == _myNewVec_61_T_3[6:0] ? myVec_82 : _GEN_8699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8701 = 7'h53 == _myNewVec_61_T_3[6:0] ? myVec_83 : _GEN_8700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8702 = 7'h54 == _myNewVec_61_T_3[6:0] ? myVec_84 : _GEN_8701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8703 = 7'h55 == _myNewVec_61_T_3[6:0] ? myVec_85 : _GEN_8702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8704 = 7'h56 == _myNewVec_61_T_3[6:0] ? myVec_86 : _GEN_8703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8705 = 7'h57 == _myNewVec_61_T_3[6:0] ? myVec_87 : _GEN_8704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8706 = 7'h58 == _myNewVec_61_T_3[6:0] ? myVec_88 : _GEN_8705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8707 = 7'h59 == _myNewVec_61_T_3[6:0] ? myVec_89 : _GEN_8706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8708 = 7'h5a == _myNewVec_61_T_3[6:0] ? myVec_90 : _GEN_8707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8709 = 7'h5b == _myNewVec_61_T_3[6:0] ? myVec_91 : _GEN_8708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8710 = 7'h5c == _myNewVec_61_T_3[6:0] ? myVec_92 : _GEN_8709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8711 = 7'h5d == _myNewVec_61_T_3[6:0] ? myVec_93 : _GEN_8710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8712 = 7'h5e == _myNewVec_61_T_3[6:0] ? myVec_94 : _GEN_8711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8713 = 7'h5f == _myNewVec_61_T_3[6:0] ? myVec_95 : _GEN_8712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8714 = 7'h60 == _myNewVec_61_T_3[6:0] ? myVec_96 : _GEN_8713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8715 = 7'h61 == _myNewVec_61_T_3[6:0] ? myVec_97 : _GEN_8714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8716 = 7'h62 == _myNewVec_61_T_3[6:0] ? myVec_98 : _GEN_8715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8717 = 7'h63 == _myNewVec_61_T_3[6:0] ? myVec_99 : _GEN_8716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8718 = 7'h64 == _myNewVec_61_T_3[6:0] ? myVec_100 : _GEN_8717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8719 = 7'h65 == _myNewVec_61_T_3[6:0] ? myVec_101 : _GEN_8718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8720 = 7'h66 == _myNewVec_61_T_3[6:0] ? myVec_102 : _GEN_8719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8721 = 7'h67 == _myNewVec_61_T_3[6:0] ? myVec_103 : _GEN_8720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8722 = 7'h68 == _myNewVec_61_T_3[6:0] ? myVec_104 : _GEN_8721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8723 = 7'h69 == _myNewVec_61_T_3[6:0] ? myVec_105 : _GEN_8722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8724 = 7'h6a == _myNewVec_61_T_3[6:0] ? myVec_106 : _GEN_8723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8725 = 7'h6b == _myNewVec_61_T_3[6:0] ? myVec_107 : _GEN_8724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8726 = 7'h6c == _myNewVec_61_T_3[6:0] ? myVec_108 : _GEN_8725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8727 = 7'h6d == _myNewVec_61_T_3[6:0] ? myVec_109 : _GEN_8726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8728 = 7'h6e == _myNewVec_61_T_3[6:0] ? myVec_110 : _GEN_8727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8729 = 7'h6f == _myNewVec_61_T_3[6:0] ? myVec_111 : _GEN_8728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8730 = 7'h70 == _myNewVec_61_T_3[6:0] ? myVec_112 : _GEN_8729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8731 = 7'h71 == _myNewVec_61_T_3[6:0] ? myVec_113 : _GEN_8730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8732 = 7'h72 == _myNewVec_61_T_3[6:0] ? myVec_114 : _GEN_8731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8733 = 7'h73 == _myNewVec_61_T_3[6:0] ? myVec_115 : _GEN_8732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8734 = 7'h74 == _myNewVec_61_T_3[6:0] ? myVec_116 : _GEN_8733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8735 = 7'h75 == _myNewVec_61_T_3[6:0] ? myVec_117 : _GEN_8734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8736 = 7'h76 == _myNewVec_61_T_3[6:0] ? myVec_118 : _GEN_8735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8737 = 7'h77 == _myNewVec_61_T_3[6:0] ? myVec_119 : _GEN_8736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8738 = 7'h78 == _myNewVec_61_T_3[6:0] ? myVec_120 : _GEN_8737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8739 = 7'h79 == _myNewVec_61_T_3[6:0] ? myVec_121 : _GEN_8738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8740 = 7'h7a == _myNewVec_61_T_3[6:0] ? myVec_122 : _GEN_8739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8741 = 7'h7b == _myNewVec_61_T_3[6:0] ? myVec_123 : _GEN_8740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8742 = 7'h7c == _myNewVec_61_T_3[6:0] ? myVec_124 : _GEN_8741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8743 = 7'h7d == _myNewVec_61_T_3[6:0] ? myVec_125 : _GEN_8742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8744 = 7'h7e == _myNewVec_61_T_3[6:0] ? myVec_126 : _GEN_8743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_61 = 7'h7f == _myNewVec_61_T_3[6:0] ? myVec_127 : _GEN_8744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_60_T_3 = _myNewVec_127_T_1 + 16'h43; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_8747 = 7'h1 == _myNewVec_60_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8748 = 7'h2 == _myNewVec_60_T_3[6:0] ? myVec_2 : _GEN_8747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8749 = 7'h3 == _myNewVec_60_T_3[6:0] ? myVec_3 : _GEN_8748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8750 = 7'h4 == _myNewVec_60_T_3[6:0] ? myVec_4 : _GEN_8749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8751 = 7'h5 == _myNewVec_60_T_3[6:0] ? myVec_5 : _GEN_8750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8752 = 7'h6 == _myNewVec_60_T_3[6:0] ? myVec_6 : _GEN_8751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8753 = 7'h7 == _myNewVec_60_T_3[6:0] ? myVec_7 : _GEN_8752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8754 = 7'h8 == _myNewVec_60_T_3[6:0] ? myVec_8 : _GEN_8753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8755 = 7'h9 == _myNewVec_60_T_3[6:0] ? myVec_9 : _GEN_8754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8756 = 7'ha == _myNewVec_60_T_3[6:0] ? myVec_10 : _GEN_8755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8757 = 7'hb == _myNewVec_60_T_3[6:0] ? myVec_11 : _GEN_8756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8758 = 7'hc == _myNewVec_60_T_3[6:0] ? myVec_12 : _GEN_8757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8759 = 7'hd == _myNewVec_60_T_3[6:0] ? myVec_13 : _GEN_8758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8760 = 7'he == _myNewVec_60_T_3[6:0] ? myVec_14 : _GEN_8759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8761 = 7'hf == _myNewVec_60_T_3[6:0] ? myVec_15 : _GEN_8760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8762 = 7'h10 == _myNewVec_60_T_3[6:0] ? myVec_16 : _GEN_8761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8763 = 7'h11 == _myNewVec_60_T_3[6:0] ? myVec_17 : _GEN_8762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8764 = 7'h12 == _myNewVec_60_T_3[6:0] ? myVec_18 : _GEN_8763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8765 = 7'h13 == _myNewVec_60_T_3[6:0] ? myVec_19 : _GEN_8764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8766 = 7'h14 == _myNewVec_60_T_3[6:0] ? myVec_20 : _GEN_8765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8767 = 7'h15 == _myNewVec_60_T_3[6:0] ? myVec_21 : _GEN_8766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8768 = 7'h16 == _myNewVec_60_T_3[6:0] ? myVec_22 : _GEN_8767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8769 = 7'h17 == _myNewVec_60_T_3[6:0] ? myVec_23 : _GEN_8768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8770 = 7'h18 == _myNewVec_60_T_3[6:0] ? myVec_24 : _GEN_8769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8771 = 7'h19 == _myNewVec_60_T_3[6:0] ? myVec_25 : _GEN_8770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8772 = 7'h1a == _myNewVec_60_T_3[6:0] ? myVec_26 : _GEN_8771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8773 = 7'h1b == _myNewVec_60_T_3[6:0] ? myVec_27 : _GEN_8772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8774 = 7'h1c == _myNewVec_60_T_3[6:0] ? myVec_28 : _GEN_8773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8775 = 7'h1d == _myNewVec_60_T_3[6:0] ? myVec_29 : _GEN_8774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8776 = 7'h1e == _myNewVec_60_T_3[6:0] ? myVec_30 : _GEN_8775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8777 = 7'h1f == _myNewVec_60_T_3[6:0] ? myVec_31 : _GEN_8776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8778 = 7'h20 == _myNewVec_60_T_3[6:0] ? myVec_32 : _GEN_8777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8779 = 7'h21 == _myNewVec_60_T_3[6:0] ? myVec_33 : _GEN_8778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8780 = 7'h22 == _myNewVec_60_T_3[6:0] ? myVec_34 : _GEN_8779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8781 = 7'h23 == _myNewVec_60_T_3[6:0] ? myVec_35 : _GEN_8780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8782 = 7'h24 == _myNewVec_60_T_3[6:0] ? myVec_36 : _GEN_8781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8783 = 7'h25 == _myNewVec_60_T_3[6:0] ? myVec_37 : _GEN_8782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8784 = 7'h26 == _myNewVec_60_T_3[6:0] ? myVec_38 : _GEN_8783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8785 = 7'h27 == _myNewVec_60_T_3[6:0] ? myVec_39 : _GEN_8784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8786 = 7'h28 == _myNewVec_60_T_3[6:0] ? myVec_40 : _GEN_8785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8787 = 7'h29 == _myNewVec_60_T_3[6:0] ? myVec_41 : _GEN_8786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8788 = 7'h2a == _myNewVec_60_T_3[6:0] ? myVec_42 : _GEN_8787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8789 = 7'h2b == _myNewVec_60_T_3[6:0] ? myVec_43 : _GEN_8788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8790 = 7'h2c == _myNewVec_60_T_3[6:0] ? myVec_44 : _GEN_8789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8791 = 7'h2d == _myNewVec_60_T_3[6:0] ? myVec_45 : _GEN_8790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8792 = 7'h2e == _myNewVec_60_T_3[6:0] ? myVec_46 : _GEN_8791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8793 = 7'h2f == _myNewVec_60_T_3[6:0] ? myVec_47 : _GEN_8792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8794 = 7'h30 == _myNewVec_60_T_3[6:0] ? myVec_48 : _GEN_8793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8795 = 7'h31 == _myNewVec_60_T_3[6:0] ? myVec_49 : _GEN_8794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8796 = 7'h32 == _myNewVec_60_T_3[6:0] ? myVec_50 : _GEN_8795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8797 = 7'h33 == _myNewVec_60_T_3[6:0] ? myVec_51 : _GEN_8796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8798 = 7'h34 == _myNewVec_60_T_3[6:0] ? myVec_52 : _GEN_8797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8799 = 7'h35 == _myNewVec_60_T_3[6:0] ? myVec_53 : _GEN_8798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8800 = 7'h36 == _myNewVec_60_T_3[6:0] ? myVec_54 : _GEN_8799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8801 = 7'h37 == _myNewVec_60_T_3[6:0] ? myVec_55 : _GEN_8800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8802 = 7'h38 == _myNewVec_60_T_3[6:0] ? myVec_56 : _GEN_8801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8803 = 7'h39 == _myNewVec_60_T_3[6:0] ? myVec_57 : _GEN_8802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8804 = 7'h3a == _myNewVec_60_T_3[6:0] ? myVec_58 : _GEN_8803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8805 = 7'h3b == _myNewVec_60_T_3[6:0] ? myVec_59 : _GEN_8804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8806 = 7'h3c == _myNewVec_60_T_3[6:0] ? myVec_60 : _GEN_8805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8807 = 7'h3d == _myNewVec_60_T_3[6:0] ? myVec_61 : _GEN_8806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8808 = 7'h3e == _myNewVec_60_T_3[6:0] ? myVec_62 : _GEN_8807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8809 = 7'h3f == _myNewVec_60_T_3[6:0] ? myVec_63 : _GEN_8808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8810 = 7'h40 == _myNewVec_60_T_3[6:0] ? myVec_64 : _GEN_8809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8811 = 7'h41 == _myNewVec_60_T_3[6:0] ? myVec_65 : _GEN_8810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8812 = 7'h42 == _myNewVec_60_T_3[6:0] ? myVec_66 : _GEN_8811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8813 = 7'h43 == _myNewVec_60_T_3[6:0] ? myVec_67 : _GEN_8812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8814 = 7'h44 == _myNewVec_60_T_3[6:0] ? myVec_68 : _GEN_8813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8815 = 7'h45 == _myNewVec_60_T_3[6:0] ? myVec_69 : _GEN_8814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8816 = 7'h46 == _myNewVec_60_T_3[6:0] ? myVec_70 : _GEN_8815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8817 = 7'h47 == _myNewVec_60_T_3[6:0] ? myVec_71 : _GEN_8816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8818 = 7'h48 == _myNewVec_60_T_3[6:0] ? myVec_72 : _GEN_8817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8819 = 7'h49 == _myNewVec_60_T_3[6:0] ? myVec_73 : _GEN_8818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8820 = 7'h4a == _myNewVec_60_T_3[6:0] ? myVec_74 : _GEN_8819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8821 = 7'h4b == _myNewVec_60_T_3[6:0] ? myVec_75 : _GEN_8820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8822 = 7'h4c == _myNewVec_60_T_3[6:0] ? myVec_76 : _GEN_8821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8823 = 7'h4d == _myNewVec_60_T_3[6:0] ? myVec_77 : _GEN_8822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8824 = 7'h4e == _myNewVec_60_T_3[6:0] ? myVec_78 : _GEN_8823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8825 = 7'h4f == _myNewVec_60_T_3[6:0] ? myVec_79 : _GEN_8824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8826 = 7'h50 == _myNewVec_60_T_3[6:0] ? myVec_80 : _GEN_8825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8827 = 7'h51 == _myNewVec_60_T_3[6:0] ? myVec_81 : _GEN_8826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8828 = 7'h52 == _myNewVec_60_T_3[6:0] ? myVec_82 : _GEN_8827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8829 = 7'h53 == _myNewVec_60_T_3[6:0] ? myVec_83 : _GEN_8828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8830 = 7'h54 == _myNewVec_60_T_3[6:0] ? myVec_84 : _GEN_8829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8831 = 7'h55 == _myNewVec_60_T_3[6:0] ? myVec_85 : _GEN_8830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8832 = 7'h56 == _myNewVec_60_T_3[6:0] ? myVec_86 : _GEN_8831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8833 = 7'h57 == _myNewVec_60_T_3[6:0] ? myVec_87 : _GEN_8832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8834 = 7'h58 == _myNewVec_60_T_3[6:0] ? myVec_88 : _GEN_8833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8835 = 7'h59 == _myNewVec_60_T_3[6:0] ? myVec_89 : _GEN_8834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8836 = 7'h5a == _myNewVec_60_T_3[6:0] ? myVec_90 : _GEN_8835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8837 = 7'h5b == _myNewVec_60_T_3[6:0] ? myVec_91 : _GEN_8836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8838 = 7'h5c == _myNewVec_60_T_3[6:0] ? myVec_92 : _GEN_8837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8839 = 7'h5d == _myNewVec_60_T_3[6:0] ? myVec_93 : _GEN_8838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8840 = 7'h5e == _myNewVec_60_T_3[6:0] ? myVec_94 : _GEN_8839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8841 = 7'h5f == _myNewVec_60_T_3[6:0] ? myVec_95 : _GEN_8840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8842 = 7'h60 == _myNewVec_60_T_3[6:0] ? myVec_96 : _GEN_8841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8843 = 7'h61 == _myNewVec_60_T_3[6:0] ? myVec_97 : _GEN_8842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8844 = 7'h62 == _myNewVec_60_T_3[6:0] ? myVec_98 : _GEN_8843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8845 = 7'h63 == _myNewVec_60_T_3[6:0] ? myVec_99 : _GEN_8844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8846 = 7'h64 == _myNewVec_60_T_3[6:0] ? myVec_100 : _GEN_8845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8847 = 7'h65 == _myNewVec_60_T_3[6:0] ? myVec_101 : _GEN_8846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8848 = 7'h66 == _myNewVec_60_T_3[6:0] ? myVec_102 : _GEN_8847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8849 = 7'h67 == _myNewVec_60_T_3[6:0] ? myVec_103 : _GEN_8848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8850 = 7'h68 == _myNewVec_60_T_3[6:0] ? myVec_104 : _GEN_8849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8851 = 7'h69 == _myNewVec_60_T_3[6:0] ? myVec_105 : _GEN_8850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8852 = 7'h6a == _myNewVec_60_T_3[6:0] ? myVec_106 : _GEN_8851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8853 = 7'h6b == _myNewVec_60_T_3[6:0] ? myVec_107 : _GEN_8852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8854 = 7'h6c == _myNewVec_60_T_3[6:0] ? myVec_108 : _GEN_8853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8855 = 7'h6d == _myNewVec_60_T_3[6:0] ? myVec_109 : _GEN_8854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8856 = 7'h6e == _myNewVec_60_T_3[6:0] ? myVec_110 : _GEN_8855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8857 = 7'h6f == _myNewVec_60_T_3[6:0] ? myVec_111 : _GEN_8856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8858 = 7'h70 == _myNewVec_60_T_3[6:0] ? myVec_112 : _GEN_8857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8859 = 7'h71 == _myNewVec_60_T_3[6:0] ? myVec_113 : _GEN_8858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8860 = 7'h72 == _myNewVec_60_T_3[6:0] ? myVec_114 : _GEN_8859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8861 = 7'h73 == _myNewVec_60_T_3[6:0] ? myVec_115 : _GEN_8860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8862 = 7'h74 == _myNewVec_60_T_3[6:0] ? myVec_116 : _GEN_8861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8863 = 7'h75 == _myNewVec_60_T_3[6:0] ? myVec_117 : _GEN_8862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8864 = 7'h76 == _myNewVec_60_T_3[6:0] ? myVec_118 : _GEN_8863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8865 = 7'h77 == _myNewVec_60_T_3[6:0] ? myVec_119 : _GEN_8864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8866 = 7'h78 == _myNewVec_60_T_3[6:0] ? myVec_120 : _GEN_8865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8867 = 7'h79 == _myNewVec_60_T_3[6:0] ? myVec_121 : _GEN_8866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8868 = 7'h7a == _myNewVec_60_T_3[6:0] ? myVec_122 : _GEN_8867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8869 = 7'h7b == _myNewVec_60_T_3[6:0] ? myVec_123 : _GEN_8868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8870 = 7'h7c == _myNewVec_60_T_3[6:0] ? myVec_124 : _GEN_8869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8871 = 7'h7d == _myNewVec_60_T_3[6:0] ? myVec_125 : _GEN_8870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8872 = 7'h7e == _myNewVec_60_T_3[6:0] ? myVec_126 : _GEN_8871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_60 = 7'h7f == _myNewVec_60_T_3[6:0] ? myVec_127 : _GEN_8872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_59_T_3 = _myNewVec_127_T_1 + 16'h44; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_8875 = 7'h1 == _myNewVec_59_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8876 = 7'h2 == _myNewVec_59_T_3[6:0] ? myVec_2 : _GEN_8875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8877 = 7'h3 == _myNewVec_59_T_3[6:0] ? myVec_3 : _GEN_8876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8878 = 7'h4 == _myNewVec_59_T_3[6:0] ? myVec_4 : _GEN_8877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8879 = 7'h5 == _myNewVec_59_T_3[6:0] ? myVec_5 : _GEN_8878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8880 = 7'h6 == _myNewVec_59_T_3[6:0] ? myVec_6 : _GEN_8879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8881 = 7'h7 == _myNewVec_59_T_3[6:0] ? myVec_7 : _GEN_8880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8882 = 7'h8 == _myNewVec_59_T_3[6:0] ? myVec_8 : _GEN_8881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8883 = 7'h9 == _myNewVec_59_T_3[6:0] ? myVec_9 : _GEN_8882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8884 = 7'ha == _myNewVec_59_T_3[6:0] ? myVec_10 : _GEN_8883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8885 = 7'hb == _myNewVec_59_T_3[6:0] ? myVec_11 : _GEN_8884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8886 = 7'hc == _myNewVec_59_T_3[6:0] ? myVec_12 : _GEN_8885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8887 = 7'hd == _myNewVec_59_T_3[6:0] ? myVec_13 : _GEN_8886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8888 = 7'he == _myNewVec_59_T_3[6:0] ? myVec_14 : _GEN_8887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8889 = 7'hf == _myNewVec_59_T_3[6:0] ? myVec_15 : _GEN_8888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8890 = 7'h10 == _myNewVec_59_T_3[6:0] ? myVec_16 : _GEN_8889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8891 = 7'h11 == _myNewVec_59_T_3[6:0] ? myVec_17 : _GEN_8890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8892 = 7'h12 == _myNewVec_59_T_3[6:0] ? myVec_18 : _GEN_8891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8893 = 7'h13 == _myNewVec_59_T_3[6:0] ? myVec_19 : _GEN_8892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8894 = 7'h14 == _myNewVec_59_T_3[6:0] ? myVec_20 : _GEN_8893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8895 = 7'h15 == _myNewVec_59_T_3[6:0] ? myVec_21 : _GEN_8894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8896 = 7'h16 == _myNewVec_59_T_3[6:0] ? myVec_22 : _GEN_8895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8897 = 7'h17 == _myNewVec_59_T_3[6:0] ? myVec_23 : _GEN_8896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8898 = 7'h18 == _myNewVec_59_T_3[6:0] ? myVec_24 : _GEN_8897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8899 = 7'h19 == _myNewVec_59_T_3[6:0] ? myVec_25 : _GEN_8898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8900 = 7'h1a == _myNewVec_59_T_3[6:0] ? myVec_26 : _GEN_8899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8901 = 7'h1b == _myNewVec_59_T_3[6:0] ? myVec_27 : _GEN_8900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8902 = 7'h1c == _myNewVec_59_T_3[6:0] ? myVec_28 : _GEN_8901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8903 = 7'h1d == _myNewVec_59_T_3[6:0] ? myVec_29 : _GEN_8902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8904 = 7'h1e == _myNewVec_59_T_3[6:0] ? myVec_30 : _GEN_8903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8905 = 7'h1f == _myNewVec_59_T_3[6:0] ? myVec_31 : _GEN_8904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8906 = 7'h20 == _myNewVec_59_T_3[6:0] ? myVec_32 : _GEN_8905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8907 = 7'h21 == _myNewVec_59_T_3[6:0] ? myVec_33 : _GEN_8906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8908 = 7'h22 == _myNewVec_59_T_3[6:0] ? myVec_34 : _GEN_8907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8909 = 7'h23 == _myNewVec_59_T_3[6:0] ? myVec_35 : _GEN_8908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8910 = 7'h24 == _myNewVec_59_T_3[6:0] ? myVec_36 : _GEN_8909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8911 = 7'h25 == _myNewVec_59_T_3[6:0] ? myVec_37 : _GEN_8910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8912 = 7'h26 == _myNewVec_59_T_3[6:0] ? myVec_38 : _GEN_8911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8913 = 7'h27 == _myNewVec_59_T_3[6:0] ? myVec_39 : _GEN_8912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8914 = 7'h28 == _myNewVec_59_T_3[6:0] ? myVec_40 : _GEN_8913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8915 = 7'h29 == _myNewVec_59_T_3[6:0] ? myVec_41 : _GEN_8914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8916 = 7'h2a == _myNewVec_59_T_3[6:0] ? myVec_42 : _GEN_8915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8917 = 7'h2b == _myNewVec_59_T_3[6:0] ? myVec_43 : _GEN_8916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8918 = 7'h2c == _myNewVec_59_T_3[6:0] ? myVec_44 : _GEN_8917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8919 = 7'h2d == _myNewVec_59_T_3[6:0] ? myVec_45 : _GEN_8918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8920 = 7'h2e == _myNewVec_59_T_3[6:0] ? myVec_46 : _GEN_8919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8921 = 7'h2f == _myNewVec_59_T_3[6:0] ? myVec_47 : _GEN_8920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8922 = 7'h30 == _myNewVec_59_T_3[6:0] ? myVec_48 : _GEN_8921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8923 = 7'h31 == _myNewVec_59_T_3[6:0] ? myVec_49 : _GEN_8922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8924 = 7'h32 == _myNewVec_59_T_3[6:0] ? myVec_50 : _GEN_8923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8925 = 7'h33 == _myNewVec_59_T_3[6:0] ? myVec_51 : _GEN_8924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8926 = 7'h34 == _myNewVec_59_T_3[6:0] ? myVec_52 : _GEN_8925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8927 = 7'h35 == _myNewVec_59_T_3[6:0] ? myVec_53 : _GEN_8926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8928 = 7'h36 == _myNewVec_59_T_3[6:0] ? myVec_54 : _GEN_8927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8929 = 7'h37 == _myNewVec_59_T_3[6:0] ? myVec_55 : _GEN_8928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8930 = 7'h38 == _myNewVec_59_T_3[6:0] ? myVec_56 : _GEN_8929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8931 = 7'h39 == _myNewVec_59_T_3[6:0] ? myVec_57 : _GEN_8930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8932 = 7'h3a == _myNewVec_59_T_3[6:0] ? myVec_58 : _GEN_8931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8933 = 7'h3b == _myNewVec_59_T_3[6:0] ? myVec_59 : _GEN_8932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8934 = 7'h3c == _myNewVec_59_T_3[6:0] ? myVec_60 : _GEN_8933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8935 = 7'h3d == _myNewVec_59_T_3[6:0] ? myVec_61 : _GEN_8934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8936 = 7'h3e == _myNewVec_59_T_3[6:0] ? myVec_62 : _GEN_8935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8937 = 7'h3f == _myNewVec_59_T_3[6:0] ? myVec_63 : _GEN_8936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8938 = 7'h40 == _myNewVec_59_T_3[6:0] ? myVec_64 : _GEN_8937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8939 = 7'h41 == _myNewVec_59_T_3[6:0] ? myVec_65 : _GEN_8938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8940 = 7'h42 == _myNewVec_59_T_3[6:0] ? myVec_66 : _GEN_8939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8941 = 7'h43 == _myNewVec_59_T_3[6:0] ? myVec_67 : _GEN_8940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8942 = 7'h44 == _myNewVec_59_T_3[6:0] ? myVec_68 : _GEN_8941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8943 = 7'h45 == _myNewVec_59_T_3[6:0] ? myVec_69 : _GEN_8942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8944 = 7'h46 == _myNewVec_59_T_3[6:0] ? myVec_70 : _GEN_8943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8945 = 7'h47 == _myNewVec_59_T_3[6:0] ? myVec_71 : _GEN_8944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8946 = 7'h48 == _myNewVec_59_T_3[6:0] ? myVec_72 : _GEN_8945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8947 = 7'h49 == _myNewVec_59_T_3[6:0] ? myVec_73 : _GEN_8946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8948 = 7'h4a == _myNewVec_59_T_3[6:0] ? myVec_74 : _GEN_8947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8949 = 7'h4b == _myNewVec_59_T_3[6:0] ? myVec_75 : _GEN_8948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8950 = 7'h4c == _myNewVec_59_T_3[6:0] ? myVec_76 : _GEN_8949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8951 = 7'h4d == _myNewVec_59_T_3[6:0] ? myVec_77 : _GEN_8950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8952 = 7'h4e == _myNewVec_59_T_3[6:0] ? myVec_78 : _GEN_8951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8953 = 7'h4f == _myNewVec_59_T_3[6:0] ? myVec_79 : _GEN_8952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8954 = 7'h50 == _myNewVec_59_T_3[6:0] ? myVec_80 : _GEN_8953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8955 = 7'h51 == _myNewVec_59_T_3[6:0] ? myVec_81 : _GEN_8954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8956 = 7'h52 == _myNewVec_59_T_3[6:0] ? myVec_82 : _GEN_8955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8957 = 7'h53 == _myNewVec_59_T_3[6:0] ? myVec_83 : _GEN_8956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8958 = 7'h54 == _myNewVec_59_T_3[6:0] ? myVec_84 : _GEN_8957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8959 = 7'h55 == _myNewVec_59_T_3[6:0] ? myVec_85 : _GEN_8958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8960 = 7'h56 == _myNewVec_59_T_3[6:0] ? myVec_86 : _GEN_8959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8961 = 7'h57 == _myNewVec_59_T_3[6:0] ? myVec_87 : _GEN_8960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8962 = 7'h58 == _myNewVec_59_T_3[6:0] ? myVec_88 : _GEN_8961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8963 = 7'h59 == _myNewVec_59_T_3[6:0] ? myVec_89 : _GEN_8962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8964 = 7'h5a == _myNewVec_59_T_3[6:0] ? myVec_90 : _GEN_8963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8965 = 7'h5b == _myNewVec_59_T_3[6:0] ? myVec_91 : _GEN_8964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8966 = 7'h5c == _myNewVec_59_T_3[6:0] ? myVec_92 : _GEN_8965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8967 = 7'h5d == _myNewVec_59_T_3[6:0] ? myVec_93 : _GEN_8966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8968 = 7'h5e == _myNewVec_59_T_3[6:0] ? myVec_94 : _GEN_8967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8969 = 7'h5f == _myNewVec_59_T_3[6:0] ? myVec_95 : _GEN_8968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8970 = 7'h60 == _myNewVec_59_T_3[6:0] ? myVec_96 : _GEN_8969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8971 = 7'h61 == _myNewVec_59_T_3[6:0] ? myVec_97 : _GEN_8970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8972 = 7'h62 == _myNewVec_59_T_3[6:0] ? myVec_98 : _GEN_8971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8973 = 7'h63 == _myNewVec_59_T_3[6:0] ? myVec_99 : _GEN_8972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8974 = 7'h64 == _myNewVec_59_T_3[6:0] ? myVec_100 : _GEN_8973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8975 = 7'h65 == _myNewVec_59_T_3[6:0] ? myVec_101 : _GEN_8974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8976 = 7'h66 == _myNewVec_59_T_3[6:0] ? myVec_102 : _GEN_8975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8977 = 7'h67 == _myNewVec_59_T_3[6:0] ? myVec_103 : _GEN_8976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8978 = 7'h68 == _myNewVec_59_T_3[6:0] ? myVec_104 : _GEN_8977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8979 = 7'h69 == _myNewVec_59_T_3[6:0] ? myVec_105 : _GEN_8978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8980 = 7'h6a == _myNewVec_59_T_3[6:0] ? myVec_106 : _GEN_8979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8981 = 7'h6b == _myNewVec_59_T_3[6:0] ? myVec_107 : _GEN_8980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8982 = 7'h6c == _myNewVec_59_T_3[6:0] ? myVec_108 : _GEN_8981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8983 = 7'h6d == _myNewVec_59_T_3[6:0] ? myVec_109 : _GEN_8982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8984 = 7'h6e == _myNewVec_59_T_3[6:0] ? myVec_110 : _GEN_8983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8985 = 7'h6f == _myNewVec_59_T_3[6:0] ? myVec_111 : _GEN_8984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8986 = 7'h70 == _myNewVec_59_T_3[6:0] ? myVec_112 : _GEN_8985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8987 = 7'h71 == _myNewVec_59_T_3[6:0] ? myVec_113 : _GEN_8986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8988 = 7'h72 == _myNewVec_59_T_3[6:0] ? myVec_114 : _GEN_8987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8989 = 7'h73 == _myNewVec_59_T_3[6:0] ? myVec_115 : _GEN_8988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8990 = 7'h74 == _myNewVec_59_T_3[6:0] ? myVec_116 : _GEN_8989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8991 = 7'h75 == _myNewVec_59_T_3[6:0] ? myVec_117 : _GEN_8990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8992 = 7'h76 == _myNewVec_59_T_3[6:0] ? myVec_118 : _GEN_8991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8993 = 7'h77 == _myNewVec_59_T_3[6:0] ? myVec_119 : _GEN_8992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8994 = 7'h78 == _myNewVec_59_T_3[6:0] ? myVec_120 : _GEN_8993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8995 = 7'h79 == _myNewVec_59_T_3[6:0] ? myVec_121 : _GEN_8994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8996 = 7'h7a == _myNewVec_59_T_3[6:0] ? myVec_122 : _GEN_8995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8997 = 7'h7b == _myNewVec_59_T_3[6:0] ? myVec_123 : _GEN_8996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8998 = 7'h7c == _myNewVec_59_T_3[6:0] ? myVec_124 : _GEN_8997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_8999 = 7'h7d == _myNewVec_59_T_3[6:0] ? myVec_125 : _GEN_8998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9000 = 7'h7e == _myNewVec_59_T_3[6:0] ? myVec_126 : _GEN_8999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_59 = 7'h7f == _myNewVec_59_T_3[6:0] ? myVec_127 : _GEN_9000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_58_T_3 = _myNewVec_127_T_1 + 16'h45; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_9003 = 7'h1 == _myNewVec_58_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9004 = 7'h2 == _myNewVec_58_T_3[6:0] ? myVec_2 : _GEN_9003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9005 = 7'h3 == _myNewVec_58_T_3[6:0] ? myVec_3 : _GEN_9004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9006 = 7'h4 == _myNewVec_58_T_3[6:0] ? myVec_4 : _GEN_9005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9007 = 7'h5 == _myNewVec_58_T_3[6:0] ? myVec_5 : _GEN_9006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9008 = 7'h6 == _myNewVec_58_T_3[6:0] ? myVec_6 : _GEN_9007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9009 = 7'h7 == _myNewVec_58_T_3[6:0] ? myVec_7 : _GEN_9008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9010 = 7'h8 == _myNewVec_58_T_3[6:0] ? myVec_8 : _GEN_9009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9011 = 7'h9 == _myNewVec_58_T_3[6:0] ? myVec_9 : _GEN_9010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9012 = 7'ha == _myNewVec_58_T_3[6:0] ? myVec_10 : _GEN_9011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9013 = 7'hb == _myNewVec_58_T_3[6:0] ? myVec_11 : _GEN_9012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9014 = 7'hc == _myNewVec_58_T_3[6:0] ? myVec_12 : _GEN_9013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9015 = 7'hd == _myNewVec_58_T_3[6:0] ? myVec_13 : _GEN_9014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9016 = 7'he == _myNewVec_58_T_3[6:0] ? myVec_14 : _GEN_9015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9017 = 7'hf == _myNewVec_58_T_3[6:0] ? myVec_15 : _GEN_9016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9018 = 7'h10 == _myNewVec_58_T_3[6:0] ? myVec_16 : _GEN_9017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9019 = 7'h11 == _myNewVec_58_T_3[6:0] ? myVec_17 : _GEN_9018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9020 = 7'h12 == _myNewVec_58_T_3[6:0] ? myVec_18 : _GEN_9019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9021 = 7'h13 == _myNewVec_58_T_3[6:0] ? myVec_19 : _GEN_9020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9022 = 7'h14 == _myNewVec_58_T_3[6:0] ? myVec_20 : _GEN_9021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9023 = 7'h15 == _myNewVec_58_T_3[6:0] ? myVec_21 : _GEN_9022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9024 = 7'h16 == _myNewVec_58_T_3[6:0] ? myVec_22 : _GEN_9023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9025 = 7'h17 == _myNewVec_58_T_3[6:0] ? myVec_23 : _GEN_9024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9026 = 7'h18 == _myNewVec_58_T_3[6:0] ? myVec_24 : _GEN_9025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9027 = 7'h19 == _myNewVec_58_T_3[6:0] ? myVec_25 : _GEN_9026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9028 = 7'h1a == _myNewVec_58_T_3[6:0] ? myVec_26 : _GEN_9027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9029 = 7'h1b == _myNewVec_58_T_3[6:0] ? myVec_27 : _GEN_9028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9030 = 7'h1c == _myNewVec_58_T_3[6:0] ? myVec_28 : _GEN_9029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9031 = 7'h1d == _myNewVec_58_T_3[6:0] ? myVec_29 : _GEN_9030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9032 = 7'h1e == _myNewVec_58_T_3[6:0] ? myVec_30 : _GEN_9031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9033 = 7'h1f == _myNewVec_58_T_3[6:0] ? myVec_31 : _GEN_9032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9034 = 7'h20 == _myNewVec_58_T_3[6:0] ? myVec_32 : _GEN_9033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9035 = 7'h21 == _myNewVec_58_T_3[6:0] ? myVec_33 : _GEN_9034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9036 = 7'h22 == _myNewVec_58_T_3[6:0] ? myVec_34 : _GEN_9035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9037 = 7'h23 == _myNewVec_58_T_3[6:0] ? myVec_35 : _GEN_9036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9038 = 7'h24 == _myNewVec_58_T_3[6:0] ? myVec_36 : _GEN_9037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9039 = 7'h25 == _myNewVec_58_T_3[6:0] ? myVec_37 : _GEN_9038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9040 = 7'h26 == _myNewVec_58_T_3[6:0] ? myVec_38 : _GEN_9039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9041 = 7'h27 == _myNewVec_58_T_3[6:0] ? myVec_39 : _GEN_9040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9042 = 7'h28 == _myNewVec_58_T_3[6:0] ? myVec_40 : _GEN_9041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9043 = 7'h29 == _myNewVec_58_T_3[6:0] ? myVec_41 : _GEN_9042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9044 = 7'h2a == _myNewVec_58_T_3[6:0] ? myVec_42 : _GEN_9043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9045 = 7'h2b == _myNewVec_58_T_3[6:0] ? myVec_43 : _GEN_9044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9046 = 7'h2c == _myNewVec_58_T_3[6:0] ? myVec_44 : _GEN_9045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9047 = 7'h2d == _myNewVec_58_T_3[6:0] ? myVec_45 : _GEN_9046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9048 = 7'h2e == _myNewVec_58_T_3[6:0] ? myVec_46 : _GEN_9047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9049 = 7'h2f == _myNewVec_58_T_3[6:0] ? myVec_47 : _GEN_9048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9050 = 7'h30 == _myNewVec_58_T_3[6:0] ? myVec_48 : _GEN_9049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9051 = 7'h31 == _myNewVec_58_T_3[6:0] ? myVec_49 : _GEN_9050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9052 = 7'h32 == _myNewVec_58_T_3[6:0] ? myVec_50 : _GEN_9051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9053 = 7'h33 == _myNewVec_58_T_3[6:0] ? myVec_51 : _GEN_9052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9054 = 7'h34 == _myNewVec_58_T_3[6:0] ? myVec_52 : _GEN_9053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9055 = 7'h35 == _myNewVec_58_T_3[6:0] ? myVec_53 : _GEN_9054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9056 = 7'h36 == _myNewVec_58_T_3[6:0] ? myVec_54 : _GEN_9055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9057 = 7'h37 == _myNewVec_58_T_3[6:0] ? myVec_55 : _GEN_9056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9058 = 7'h38 == _myNewVec_58_T_3[6:0] ? myVec_56 : _GEN_9057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9059 = 7'h39 == _myNewVec_58_T_3[6:0] ? myVec_57 : _GEN_9058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9060 = 7'h3a == _myNewVec_58_T_3[6:0] ? myVec_58 : _GEN_9059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9061 = 7'h3b == _myNewVec_58_T_3[6:0] ? myVec_59 : _GEN_9060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9062 = 7'h3c == _myNewVec_58_T_3[6:0] ? myVec_60 : _GEN_9061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9063 = 7'h3d == _myNewVec_58_T_3[6:0] ? myVec_61 : _GEN_9062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9064 = 7'h3e == _myNewVec_58_T_3[6:0] ? myVec_62 : _GEN_9063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9065 = 7'h3f == _myNewVec_58_T_3[6:0] ? myVec_63 : _GEN_9064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9066 = 7'h40 == _myNewVec_58_T_3[6:0] ? myVec_64 : _GEN_9065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9067 = 7'h41 == _myNewVec_58_T_3[6:0] ? myVec_65 : _GEN_9066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9068 = 7'h42 == _myNewVec_58_T_3[6:0] ? myVec_66 : _GEN_9067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9069 = 7'h43 == _myNewVec_58_T_3[6:0] ? myVec_67 : _GEN_9068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9070 = 7'h44 == _myNewVec_58_T_3[6:0] ? myVec_68 : _GEN_9069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9071 = 7'h45 == _myNewVec_58_T_3[6:0] ? myVec_69 : _GEN_9070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9072 = 7'h46 == _myNewVec_58_T_3[6:0] ? myVec_70 : _GEN_9071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9073 = 7'h47 == _myNewVec_58_T_3[6:0] ? myVec_71 : _GEN_9072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9074 = 7'h48 == _myNewVec_58_T_3[6:0] ? myVec_72 : _GEN_9073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9075 = 7'h49 == _myNewVec_58_T_3[6:0] ? myVec_73 : _GEN_9074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9076 = 7'h4a == _myNewVec_58_T_3[6:0] ? myVec_74 : _GEN_9075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9077 = 7'h4b == _myNewVec_58_T_3[6:0] ? myVec_75 : _GEN_9076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9078 = 7'h4c == _myNewVec_58_T_3[6:0] ? myVec_76 : _GEN_9077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9079 = 7'h4d == _myNewVec_58_T_3[6:0] ? myVec_77 : _GEN_9078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9080 = 7'h4e == _myNewVec_58_T_3[6:0] ? myVec_78 : _GEN_9079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9081 = 7'h4f == _myNewVec_58_T_3[6:0] ? myVec_79 : _GEN_9080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9082 = 7'h50 == _myNewVec_58_T_3[6:0] ? myVec_80 : _GEN_9081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9083 = 7'h51 == _myNewVec_58_T_3[6:0] ? myVec_81 : _GEN_9082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9084 = 7'h52 == _myNewVec_58_T_3[6:0] ? myVec_82 : _GEN_9083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9085 = 7'h53 == _myNewVec_58_T_3[6:0] ? myVec_83 : _GEN_9084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9086 = 7'h54 == _myNewVec_58_T_3[6:0] ? myVec_84 : _GEN_9085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9087 = 7'h55 == _myNewVec_58_T_3[6:0] ? myVec_85 : _GEN_9086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9088 = 7'h56 == _myNewVec_58_T_3[6:0] ? myVec_86 : _GEN_9087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9089 = 7'h57 == _myNewVec_58_T_3[6:0] ? myVec_87 : _GEN_9088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9090 = 7'h58 == _myNewVec_58_T_3[6:0] ? myVec_88 : _GEN_9089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9091 = 7'h59 == _myNewVec_58_T_3[6:0] ? myVec_89 : _GEN_9090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9092 = 7'h5a == _myNewVec_58_T_3[6:0] ? myVec_90 : _GEN_9091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9093 = 7'h5b == _myNewVec_58_T_3[6:0] ? myVec_91 : _GEN_9092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9094 = 7'h5c == _myNewVec_58_T_3[6:0] ? myVec_92 : _GEN_9093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9095 = 7'h5d == _myNewVec_58_T_3[6:0] ? myVec_93 : _GEN_9094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9096 = 7'h5e == _myNewVec_58_T_3[6:0] ? myVec_94 : _GEN_9095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9097 = 7'h5f == _myNewVec_58_T_3[6:0] ? myVec_95 : _GEN_9096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9098 = 7'h60 == _myNewVec_58_T_3[6:0] ? myVec_96 : _GEN_9097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9099 = 7'h61 == _myNewVec_58_T_3[6:0] ? myVec_97 : _GEN_9098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9100 = 7'h62 == _myNewVec_58_T_3[6:0] ? myVec_98 : _GEN_9099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9101 = 7'h63 == _myNewVec_58_T_3[6:0] ? myVec_99 : _GEN_9100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9102 = 7'h64 == _myNewVec_58_T_3[6:0] ? myVec_100 : _GEN_9101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9103 = 7'h65 == _myNewVec_58_T_3[6:0] ? myVec_101 : _GEN_9102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9104 = 7'h66 == _myNewVec_58_T_3[6:0] ? myVec_102 : _GEN_9103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9105 = 7'h67 == _myNewVec_58_T_3[6:0] ? myVec_103 : _GEN_9104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9106 = 7'h68 == _myNewVec_58_T_3[6:0] ? myVec_104 : _GEN_9105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9107 = 7'h69 == _myNewVec_58_T_3[6:0] ? myVec_105 : _GEN_9106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9108 = 7'h6a == _myNewVec_58_T_3[6:0] ? myVec_106 : _GEN_9107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9109 = 7'h6b == _myNewVec_58_T_3[6:0] ? myVec_107 : _GEN_9108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9110 = 7'h6c == _myNewVec_58_T_3[6:0] ? myVec_108 : _GEN_9109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9111 = 7'h6d == _myNewVec_58_T_3[6:0] ? myVec_109 : _GEN_9110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9112 = 7'h6e == _myNewVec_58_T_3[6:0] ? myVec_110 : _GEN_9111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9113 = 7'h6f == _myNewVec_58_T_3[6:0] ? myVec_111 : _GEN_9112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9114 = 7'h70 == _myNewVec_58_T_3[6:0] ? myVec_112 : _GEN_9113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9115 = 7'h71 == _myNewVec_58_T_3[6:0] ? myVec_113 : _GEN_9114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9116 = 7'h72 == _myNewVec_58_T_3[6:0] ? myVec_114 : _GEN_9115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9117 = 7'h73 == _myNewVec_58_T_3[6:0] ? myVec_115 : _GEN_9116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9118 = 7'h74 == _myNewVec_58_T_3[6:0] ? myVec_116 : _GEN_9117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9119 = 7'h75 == _myNewVec_58_T_3[6:0] ? myVec_117 : _GEN_9118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9120 = 7'h76 == _myNewVec_58_T_3[6:0] ? myVec_118 : _GEN_9119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9121 = 7'h77 == _myNewVec_58_T_3[6:0] ? myVec_119 : _GEN_9120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9122 = 7'h78 == _myNewVec_58_T_3[6:0] ? myVec_120 : _GEN_9121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9123 = 7'h79 == _myNewVec_58_T_3[6:0] ? myVec_121 : _GEN_9122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9124 = 7'h7a == _myNewVec_58_T_3[6:0] ? myVec_122 : _GEN_9123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9125 = 7'h7b == _myNewVec_58_T_3[6:0] ? myVec_123 : _GEN_9124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9126 = 7'h7c == _myNewVec_58_T_3[6:0] ? myVec_124 : _GEN_9125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9127 = 7'h7d == _myNewVec_58_T_3[6:0] ? myVec_125 : _GEN_9126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9128 = 7'h7e == _myNewVec_58_T_3[6:0] ? myVec_126 : _GEN_9127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_58 = 7'h7f == _myNewVec_58_T_3[6:0] ? myVec_127 : _GEN_9128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_57_T_3 = _myNewVec_127_T_1 + 16'h46; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_9131 = 7'h1 == _myNewVec_57_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9132 = 7'h2 == _myNewVec_57_T_3[6:0] ? myVec_2 : _GEN_9131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9133 = 7'h3 == _myNewVec_57_T_3[6:0] ? myVec_3 : _GEN_9132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9134 = 7'h4 == _myNewVec_57_T_3[6:0] ? myVec_4 : _GEN_9133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9135 = 7'h5 == _myNewVec_57_T_3[6:0] ? myVec_5 : _GEN_9134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9136 = 7'h6 == _myNewVec_57_T_3[6:0] ? myVec_6 : _GEN_9135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9137 = 7'h7 == _myNewVec_57_T_3[6:0] ? myVec_7 : _GEN_9136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9138 = 7'h8 == _myNewVec_57_T_3[6:0] ? myVec_8 : _GEN_9137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9139 = 7'h9 == _myNewVec_57_T_3[6:0] ? myVec_9 : _GEN_9138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9140 = 7'ha == _myNewVec_57_T_3[6:0] ? myVec_10 : _GEN_9139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9141 = 7'hb == _myNewVec_57_T_3[6:0] ? myVec_11 : _GEN_9140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9142 = 7'hc == _myNewVec_57_T_3[6:0] ? myVec_12 : _GEN_9141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9143 = 7'hd == _myNewVec_57_T_3[6:0] ? myVec_13 : _GEN_9142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9144 = 7'he == _myNewVec_57_T_3[6:0] ? myVec_14 : _GEN_9143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9145 = 7'hf == _myNewVec_57_T_3[6:0] ? myVec_15 : _GEN_9144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9146 = 7'h10 == _myNewVec_57_T_3[6:0] ? myVec_16 : _GEN_9145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9147 = 7'h11 == _myNewVec_57_T_3[6:0] ? myVec_17 : _GEN_9146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9148 = 7'h12 == _myNewVec_57_T_3[6:0] ? myVec_18 : _GEN_9147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9149 = 7'h13 == _myNewVec_57_T_3[6:0] ? myVec_19 : _GEN_9148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9150 = 7'h14 == _myNewVec_57_T_3[6:0] ? myVec_20 : _GEN_9149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9151 = 7'h15 == _myNewVec_57_T_3[6:0] ? myVec_21 : _GEN_9150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9152 = 7'h16 == _myNewVec_57_T_3[6:0] ? myVec_22 : _GEN_9151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9153 = 7'h17 == _myNewVec_57_T_3[6:0] ? myVec_23 : _GEN_9152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9154 = 7'h18 == _myNewVec_57_T_3[6:0] ? myVec_24 : _GEN_9153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9155 = 7'h19 == _myNewVec_57_T_3[6:0] ? myVec_25 : _GEN_9154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9156 = 7'h1a == _myNewVec_57_T_3[6:0] ? myVec_26 : _GEN_9155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9157 = 7'h1b == _myNewVec_57_T_3[6:0] ? myVec_27 : _GEN_9156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9158 = 7'h1c == _myNewVec_57_T_3[6:0] ? myVec_28 : _GEN_9157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9159 = 7'h1d == _myNewVec_57_T_3[6:0] ? myVec_29 : _GEN_9158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9160 = 7'h1e == _myNewVec_57_T_3[6:0] ? myVec_30 : _GEN_9159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9161 = 7'h1f == _myNewVec_57_T_3[6:0] ? myVec_31 : _GEN_9160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9162 = 7'h20 == _myNewVec_57_T_3[6:0] ? myVec_32 : _GEN_9161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9163 = 7'h21 == _myNewVec_57_T_3[6:0] ? myVec_33 : _GEN_9162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9164 = 7'h22 == _myNewVec_57_T_3[6:0] ? myVec_34 : _GEN_9163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9165 = 7'h23 == _myNewVec_57_T_3[6:0] ? myVec_35 : _GEN_9164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9166 = 7'h24 == _myNewVec_57_T_3[6:0] ? myVec_36 : _GEN_9165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9167 = 7'h25 == _myNewVec_57_T_3[6:0] ? myVec_37 : _GEN_9166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9168 = 7'h26 == _myNewVec_57_T_3[6:0] ? myVec_38 : _GEN_9167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9169 = 7'h27 == _myNewVec_57_T_3[6:0] ? myVec_39 : _GEN_9168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9170 = 7'h28 == _myNewVec_57_T_3[6:0] ? myVec_40 : _GEN_9169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9171 = 7'h29 == _myNewVec_57_T_3[6:0] ? myVec_41 : _GEN_9170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9172 = 7'h2a == _myNewVec_57_T_3[6:0] ? myVec_42 : _GEN_9171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9173 = 7'h2b == _myNewVec_57_T_3[6:0] ? myVec_43 : _GEN_9172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9174 = 7'h2c == _myNewVec_57_T_3[6:0] ? myVec_44 : _GEN_9173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9175 = 7'h2d == _myNewVec_57_T_3[6:0] ? myVec_45 : _GEN_9174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9176 = 7'h2e == _myNewVec_57_T_3[6:0] ? myVec_46 : _GEN_9175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9177 = 7'h2f == _myNewVec_57_T_3[6:0] ? myVec_47 : _GEN_9176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9178 = 7'h30 == _myNewVec_57_T_3[6:0] ? myVec_48 : _GEN_9177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9179 = 7'h31 == _myNewVec_57_T_3[6:0] ? myVec_49 : _GEN_9178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9180 = 7'h32 == _myNewVec_57_T_3[6:0] ? myVec_50 : _GEN_9179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9181 = 7'h33 == _myNewVec_57_T_3[6:0] ? myVec_51 : _GEN_9180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9182 = 7'h34 == _myNewVec_57_T_3[6:0] ? myVec_52 : _GEN_9181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9183 = 7'h35 == _myNewVec_57_T_3[6:0] ? myVec_53 : _GEN_9182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9184 = 7'h36 == _myNewVec_57_T_3[6:0] ? myVec_54 : _GEN_9183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9185 = 7'h37 == _myNewVec_57_T_3[6:0] ? myVec_55 : _GEN_9184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9186 = 7'h38 == _myNewVec_57_T_3[6:0] ? myVec_56 : _GEN_9185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9187 = 7'h39 == _myNewVec_57_T_3[6:0] ? myVec_57 : _GEN_9186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9188 = 7'h3a == _myNewVec_57_T_3[6:0] ? myVec_58 : _GEN_9187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9189 = 7'h3b == _myNewVec_57_T_3[6:0] ? myVec_59 : _GEN_9188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9190 = 7'h3c == _myNewVec_57_T_3[6:0] ? myVec_60 : _GEN_9189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9191 = 7'h3d == _myNewVec_57_T_3[6:0] ? myVec_61 : _GEN_9190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9192 = 7'h3e == _myNewVec_57_T_3[6:0] ? myVec_62 : _GEN_9191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9193 = 7'h3f == _myNewVec_57_T_3[6:0] ? myVec_63 : _GEN_9192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9194 = 7'h40 == _myNewVec_57_T_3[6:0] ? myVec_64 : _GEN_9193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9195 = 7'h41 == _myNewVec_57_T_3[6:0] ? myVec_65 : _GEN_9194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9196 = 7'h42 == _myNewVec_57_T_3[6:0] ? myVec_66 : _GEN_9195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9197 = 7'h43 == _myNewVec_57_T_3[6:0] ? myVec_67 : _GEN_9196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9198 = 7'h44 == _myNewVec_57_T_3[6:0] ? myVec_68 : _GEN_9197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9199 = 7'h45 == _myNewVec_57_T_3[6:0] ? myVec_69 : _GEN_9198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9200 = 7'h46 == _myNewVec_57_T_3[6:0] ? myVec_70 : _GEN_9199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9201 = 7'h47 == _myNewVec_57_T_3[6:0] ? myVec_71 : _GEN_9200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9202 = 7'h48 == _myNewVec_57_T_3[6:0] ? myVec_72 : _GEN_9201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9203 = 7'h49 == _myNewVec_57_T_3[6:0] ? myVec_73 : _GEN_9202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9204 = 7'h4a == _myNewVec_57_T_3[6:0] ? myVec_74 : _GEN_9203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9205 = 7'h4b == _myNewVec_57_T_3[6:0] ? myVec_75 : _GEN_9204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9206 = 7'h4c == _myNewVec_57_T_3[6:0] ? myVec_76 : _GEN_9205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9207 = 7'h4d == _myNewVec_57_T_3[6:0] ? myVec_77 : _GEN_9206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9208 = 7'h4e == _myNewVec_57_T_3[6:0] ? myVec_78 : _GEN_9207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9209 = 7'h4f == _myNewVec_57_T_3[6:0] ? myVec_79 : _GEN_9208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9210 = 7'h50 == _myNewVec_57_T_3[6:0] ? myVec_80 : _GEN_9209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9211 = 7'h51 == _myNewVec_57_T_3[6:0] ? myVec_81 : _GEN_9210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9212 = 7'h52 == _myNewVec_57_T_3[6:0] ? myVec_82 : _GEN_9211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9213 = 7'h53 == _myNewVec_57_T_3[6:0] ? myVec_83 : _GEN_9212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9214 = 7'h54 == _myNewVec_57_T_3[6:0] ? myVec_84 : _GEN_9213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9215 = 7'h55 == _myNewVec_57_T_3[6:0] ? myVec_85 : _GEN_9214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9216 = 7'h56 == _myNewVec_57_T_3[6:0] ? myVec_86 : _GEN_9215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9217 = 7'h57 == _myNewVec_57_T_3[6:0] ? myVec_87 : _GEN_9216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9218 = 7'h58 == _myNewVec_57_T_3[6:0] ? myVec_88 : _GEN_9217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9219 = 7'h59 == _myNewVec_57_T_3[6:0] ? myVec_89 : _GEN_9218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9220 = 7'h5a == _myNewVec_57_T_3[6:0] ? myVec_90 : _GEN_9219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9221 = 7'h5b == _myNewVec_57_T_3[6:0] ? myVec_91 : _GEN_9220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9222 = 7'h5c == _myNewVec_57_T_3[6:0] ? myVec_92 : _GEN_9221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9223 = 7'h5d == _myNewVec_57_T_3[6:0] ? myVec_93 : _GEN_9222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9224 = 7'h5e == _myNewVec_57_T_3[6:0] ? myVec_94 : _GEN_9223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9225 = 7'h5f == _myNewVec_57_T_3[6:0] ? myVec_95 : _GEN_9224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9226 = 7'h60 == _myNewVec_57_T_3[6:0] ? myVec_96 : _GEN_9225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9227 = 7'h61 == _myNewVec_57_T_3[6:0] ? myVec_97 : _GEN_9226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9228 = 7'h62 == _myNewVec_57_T_3[6:0] ? myVec_98 : _GEN_9227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9229 = 7'h63 == _myNewVec_57_T_3[6:0] ? myVec_99 : _GEN_9228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9230 = 7'h64 == _myNewVec_57_T_3[6:0] ? myVec_100 : _GEN_9229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9231 = 7'h65 == _myNewVec_57_T_3[6:0] ? myVec_101 : _GEN_9230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9232 = 7'h66 == _myNewVec_57_T_3[6:0] ? myVec_102 : _GEN_9231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9233 = 7'h67 == _myNewVec_57_T_3[6:0] ? myVec_103 : _GEN_9232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9234 = 7'h68 == _myNewVec_57_T_3[6:0] ? myVec_104 : _GEN_9233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9235 = 7'h69 == _myNewVec_57_T_3[6:0] ? myVec_105 : _GEN_9234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9236 = 7'h6a == _myNewVec_57_T_3[6:0] ? myVec_106 : _GEN_9235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9237 = 7'h6b == _myNewVec_57_T_3[6:0] ? myVec_107 : _GEN_9236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9238 = 7'h6c == _myNewVec_57_T_3[6:0] ? myVec_108 : _GEN_9237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9239 = 7'h6d == _myNewVec_57_T_3[6:0] ? myVec_109 : _GEN_9238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9240 = 7'h6e == _myNewVec_57_T_3[6:0] ? myVec_110 : _GEN_9239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9241 = 7'h6f == _myNewVec_57_T_3[6:0] ? myVec_111 : _GEN_9240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9242 = 7'h70 == _myNewVec_57_T_3[6:0] ? myVec_112 : _GEN_9241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9243 = 7'h71 == _myNewVec_57_T_3[6:0] ? myVec_113 : _GEN_9242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9244 = 7'h72 == _myNewVec_57_T_3[6:0] ? myVec_114 : _GEN_9243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9245 = 7'h73 == _myNewVec_57_T_3[6:0] ? myVec_115 : _GEN_9244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9246 = 7'h74 == _myNewVec_57_T_3[6:0] ? myVec_116 : _GEN_9245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9247 = 7'h75 == _myNewVec_57_T_3[6:0] ? myVec_117 : _GEN_9246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9248 = 7'h76 == _myNewVec_57_T_3[6:0] ? myVec_118 : _GEN_9247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9249 = 7'h77 == _myNewVec_57_T_3[6:0] ? myVec_119 : _GEN_9248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9250 = 7'h78 == _myNewVec_57_T_3[6:0] ? myVec_120 : _GEN_9249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9251 = 7'h79 == _myNewVec_57_T_3[6:0] ? myVec_121 : _GEN_9250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9252 = 7'h7a == _myNewVec_57_T_3[6:0] ? myVec_122 : _GEN_9251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9253 = 7'h7b == _myNewVec_57_T_3[6:0] ? myVec_123 : _GEN_9252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9254 = 7'h7c == _myNewVec_57_T_3[6:0] ? myVec_124 : _GEN_9253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9255 = 7'h7d == _myNewVec_57_T_3[6:0] ? myVec_125 : _GEN_9254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9256 = 7'h7e == _myNewVec_57_T_3[6:0] ? myVec_126 : _GEN_9255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_57 = 7'h7f == _myNewVec_57_T_3[6:0] ? myVec_127 : _GEN_9256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_56_T_3 = _myNewVec_127_T_1 + 16'h47; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_9259 = 7'h1 == _myNewVec_56_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9260 = 7'h2 == _myNewVec_56_T_3[6:0] ? myVec_2 : _GEN_9259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9261 = 7'h3 == _myNewVec_56_T_3[6:0] ? myVec_3 : _GEN_9260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9262 = 7'h4 == _myNewVec_56_T_3[6:0] ? myVec_4 : _GEN_9261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9263 = 7'h5 == _myNewVec_56_T_3[6:0] ? myVec_5 : _GEN_9262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9264 = 7'h6 == _myNewVec_56_T_3[6:0] ? myVec_6 : _GEN_9263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9265 = 7'h7 == _myNewVec_56_T_3[6:0] ? myVec_7 : _GEN_9264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9266 = 7'h8 == _myNewVec_56_T_3[6:0] ? myVec_8 : _GEN_9265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9267 = 7'h9 == _myNewVec_56_T_3[6:0] ? myVec_9 : _GEN_9266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9268 = 7'ha == _myNewVec_56_T_3[6:0] ? myVec_10 : _GEN_9267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9269 = 7'hb == _myNewVec_56_T_3[6:0] ? myVec_11 : _GEN_9268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9270 = 7'hc == _myNewVec_56_T_3[6:0] ? myVec_12 : _GEN_9269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9271 = 7'hd == _myNewVec_56_T_3[6:0] ? myVec_13 : _GEN_9270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9272 = 7'he == _myNewVec_56_T_3[6:0] ? myVec_14 : _GEN_9271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9273 = 7'hf == _myNewVec_56_T_3[6:0] ? myVec_15 : _GEN_9272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9274 = 7'h10 == _myNewVec_56_T_3[6:0] ? myVec_16 : _GEN_9273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9275 = 7'h11 == _myNewVec_56_T_3[6:0] ? myVec_17 : _GEN_9274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9276 = 7'h12 == _myNewVec_56_T_3[6:0] ? myVec_18 : _GEN_9275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9277 = 7'h13 == _myNewVec_56_T_3[6:0] ? myVec_19 : _GEN_9276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9278 = 7'h14 == _myNewVec_56_T_3[6:0] ? myVec_20 : _GEN_9277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9279 = 7'h15 == _myNewVec_56_T_3[6:0] ? myVec_21 : _GEN_9278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9280 = 7'h16 == _myNewVec_56_T_3[6:0] ? myVec_22 : _GEN_9279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9281 = 7'h17 == _myNewVec_56_T_3[6:0] ? myVec_23 : _GEN_9280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9282 = 7'h18 == _myNewVec_56_T_3[6:0] ? myVec_24 : _GEN_9281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9283 = 7'h19 == _myNewVec_56_T_3[6:0] ? myVec_25 : _GEN_9282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9284 = 7'h1a == _myNewVec_56_T_3[6:0] ? myVec_26 : _GEN_9283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9285 = 7'h1b == _myNewVec_56_T_3[6:0] ? myVec_27 : _GEN_9284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9286 = 7'h1c == _myNewVec_56_T_3[6:0] ? myVec_28 : _GEN_9285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9287 = 7'h1d == _myNewVec_56_T_3[6:0] ? myVec_29 : _GEN_9286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9288 = 7'h1e == _myNewVec_56_T_3[6:0] ? myVec_30 : _GEN_9287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9289 = 7'h1f == _myNewVec_56_T_3[6:0] ? myVec_31 : _GEN_9288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9290 = 7'h20 == _myNewVec_56_T_3[6:0] ? myVec_32 : _GEN_9289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9291 = 7'h21 == _myNewVec_56_T_3[6:0] ? myVec_33 : _GEN_9290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9292 = 7'h22 == _myNewVec_56_T_3[6:0] ? myVec_34 : _GEN_9291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9293 = 7'h23 == _myNewVec_56_T_3[6:0] ? myVec_35 : _GEN_9292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9294 = 7'h24 == _myNewVec_56_T_3[6:0] ? myVec_36 : _GEN_9293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9295 = 7'h25 == _myNewVec_56_T_3[6:0] ? myVec_37 : _GEN_9294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9296 = 7'h26 == _myNewVec_56_T_3[6:0] ? myVec_38 : _GEN_9295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9297 = 7'h27 == _myNewVec_56_T_3[6:0] ? myVec_39 : _GEN_9296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9298 = 7'h28 == _myNewVec_56_T_3[6:0] ? myVec_40 : _GEN_9297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9299 = 7'h29 == _myNewVec_56_T_3[6:0] ? myVec_41 : _GEN_9298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9300 = 7'h2a == _myNewVec_56_T_3[6:0] ? myVec_42 : _GEN_9299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9301 = 7'h2b == _myNewVec_56_T_3[6:0] ? myVec_43 : _GEN_9300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9302 = 7'h2c == _myNewVec_56_T_3[6:0] ? myVec_44 : _GEN_9301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9303 = 7'h2d == _myNewVec_56_T_3[6:0] ? myVec_45 : _GEN_9302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9304 = 7'h2e == _myNewVec_56_T_3[6:0] ? myVec_46 : _GEN_9303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9305 = 7'h2f == _myNewVec_56_T_3[6:0] ? myVec_47 : _GEN_9304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9306 = 7'h30 == _myNewVec_56_T_3[6:0] ? myVec_48 : _GEN_9305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9307 = 7'h31 == _myNewVec_56_T_3[6:0] ? myVec_49 : _GEN_9306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9308 = 7'h32 == _myNewVec_56_T_3[6:0] ? myVec_50 : _GEN_9307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9309 = 7'h33 == _myNewVec_56_T_3[6:0] ? myVec_51 : _GEN_9308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9310 = 7'h34 == _myNewVec_56_T_3[6:0] ? myVec_52 : _GEN_9309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9311 = 7'h35 == _myNewVec_56_T_3[6:0] ? myVec_53 : _GEN_9310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9312 = 7'h36 == _myNewVec_56_T_3[6:0] ? myVec_54 : _GEN_9311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9313 = 7'h37 == _myNewVec_56_T_3[6:0] ? myVec_55 : _GEN_9312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9314 = 7'h38 == _myNewVec_56_T_3[6:0] ? myVec_56 : _GEN_9313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9315 = 7'h39 == _myNewVec_56_T_3[6:0] ? myVec_57 : _GEN_9314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9316 = 7'h3a == _myNewVec_56_T_3[6:0] ? myVec_58 : _GEN_9315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9317 = 7'h3b == _myNewVec_56_T_3[6:0] ? myVec_59 : _GEN_9316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9318 = 7'h3c == _myNewVec_56_T_3[6:0] ? myVec_60 : _GEN_9317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9319 = 7'h3d == _myNewVec_56_T_3[6:0] ? myVec_61 : _GEN_9318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9320 = 7'h3e == _myNewVec_56_T_3[6:0] ? myVec_62 : _GEN_9319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9321 = 7'h3f == _myNewVec_56_T_3[6:0] ? myVec_63 : _GEN_9320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9322 = 7'h40 == _myNewVec_56_T_3[6:0] ? myVec_64 : _GEN_9321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9323 = 7'h41 == _myNewVec_56_T_3[6:0] ? myVec_65 : _GEN_9322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9324 = 7'h42 == _myNewVec_56_T_3[6:0] ? myVec_66 : _GEN_9323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9325 = 7'h43 == _myNewVec_56_T_3[6:0] ? myVec_67 : _GEN_9324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9326 = 7'h44 == _myNewVec_56_T_3[6:0] ? myVec_68 : _GEN_9325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9327 = 7'h45 == _myNewVec_56_T_3[6:0] ? myVec_69 : _GEN_9326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9328 = 7'h46 == _myNewVec_56_T_3[6:0] ? myVec_70 : _GEN_9327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9329 = 7'h47 == _myNewVec_56_T_3[6:0] ? myVec_71 : _GEN_9328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9330 = 7'h48 == _myNewVec_56_T_3[6:0] ? myVec_72 : _GEN_9329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9331 = 7'h49 == _myNewVec_56_T_3[6:0] ? myVec_73 : _GEN_9330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9332 = 7'h4a == _myNewVec_56_T_3[6:0] ? myVec_74 : _GEN_9331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9333 = 7'h4b == _myNewVec_56_T_3[6:0] ? myVec_75 : _GEN_9332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9334 = 7'h4c == _myNewVec_56_T_3[6:0] ? myVec_76 : _GEN_9333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9335 = 7'h4d == _myNewVec_56_T_3[6:0] ? myVec_77 : _GEN_9334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9336 = 7'h4e == _myNewVec_56_T_3[6:0] ? myVec_78 : _GEN_9335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9337 = 7'h4f == _myNewVec_56_T_3[6:0] ? myVec_79 : _GEN_9336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9338 = 7'h50 == _myNewVec_56_T_3[6:0] ? myVec_80 : _GEN_9337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9339 = 7'h51 == _myNewVec_56_T_3[6:0] ? myVec_81 : _GEN_9338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9340 = 7'h52 == _myNewVec_56_T_3[6:0] ? myVec_82 : _GEN_9339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9341 = 7'h53 == _myNewVec_56_T_3[6:0] ? myVec_83 : _GEN_9340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9342 = 7'h54 == _myNewVec_56_T_3[6:0] ? myVec_84 : _GEN_9341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9343 = 7'h55 == _myNewVec_56_T_3[6:0] ? myVec_85 : _GEN_9342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9344 = 7'h56 == _myNewVec_56_T_3[6:0] ? myVec_86 : _GEN_9343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9345 = 7'h57 == _myNewVec_56_T_3[6:0] ? myVec_87 : _GEN_9344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9346 = 7'h58 == _myNewVec_56_T_3[6:0] ? myVec_88 : _GEN_9345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9347 = 7'h59 == _myNewVec_56_T_3[6:0] ? myVec_89 : _GEN_9346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9348 = 7'h5a == _myNewVec_56_T_3[6:0] ? myVec_90 : _GEN_9347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9349 = 7'h5b == _myNewVec_56_T_3[6:0] ? myVec_91 : _GEN_9348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9350 = 7'h5c == _myNewVec_56_T_3[6:0] ? myVec_92 : _GEN_9349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9351 = 7'h5d == _myNewVec_56_T_3[6:0] ? myVec_93 : _GEN_9350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9352 = 7'h5e == _myNewVec_56_T_3[6:0] ? myVec_94 : _GEN_9351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9353 = 7'h5f == _myNewVec_56_T_3[6:0] ? myVec_95 : _GEN_9352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9354 = 7'h60 == _myNewVec_56_T_3[6:0] ? myVec_96 : _GEN_9353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9355 = 7'h61 == _myNewVec_56_T_3[6:0] ? myVec_97 : _GEN_9354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9356 = 7'h62 == _myNewVec_56_T_3[6:0] ? myVec_98 : _GEN_9355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9357 = 7'h63 == _myNewVec_56_T_3[6:0] ? myVec_99 : _GEN_9356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9358 = 7'h64 == _myNewVec_56_T_3[6:0] ? myVec_100 : _GEN_9357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9359 = 7'h65 == _myNewVec_56_T_3[6:0] ? myVec_101 : _GEN_9358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9360 = 7'h66 == _myNewVec_56_T_3[6:0] ? myVec_102 : _GEN_9359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9361 = 7'h67 == _myNewVec_56_T_3[6:0] ? myVec_103 : _GEN_9360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9362 = 7'h68 == _myNewVec_56_T_3[6:0] ? myVec_104 : _GEN_9361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9363 = 7'h69 == _myNewVec_56_T_3[6:0] ? myVec_105 : _GEN_9362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9364 = 7'h6a == _myNewVec_56_T_3[6:0] ? myVec_106 : _GEN_9363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9365 = 7'h6b == _myNewVec_56_T_3[6:0] ? myVec_107 : _GEN_9364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9366 = 7'h6c == _myNewVec_56_T_3[6:0] ? myVec_108 : _GEN_9365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9367 = 7'h6d == _myNewVec_56_T_3[6:0] ? myVec_109 : _GEN_9366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9368 = 7'h6e == _myNewVec_56_T_3[6:0] ? myVec_110 : _GEN_9367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9369 = 7'h6f == _myNewVec_56_T_3[6:0] ? myVec_111 : _GEN_9368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9370 = 7'h70 == _myNewVec_56_T_3[6:0] ? myVec_112 : _GEN_9369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9371 = 7'h71 == _myNewVec_56_T_3[6:0] ? myVec_113 : _GEN_9370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9372 = 7'h72 == _myNewVec_56_T_3[6:0] ? myVec_114 : _GEN_9371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9373 = 7'h73 == _myNewVec_56_T_3[6:0] ? myVec_115 : _GEN_9372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9374 = 7'h74 == _myNewVec_56_T_3[6:0] ? myVec_116 : _GEN_9373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9375 = 7'h75 == _myNewVec_56_T_3[6:0] ? myVec_117 : _GEN_9374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9376 = 7'h76 == _myNewVec_56_T_3[6:0] ? myVec_118 : _GEN_9375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9377 = 7'h77 == _myNewVec_56_T_3[6:0] ? myVec_119 : _GEN_9376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9378 = 7'h78 == _myNewVec_56_T_3[6:0] ? myVec_120 : _GEN_9377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9379 = 7'h79 == _myNewVec_56_T_3[6:0] ? myVec_121 : _GEN_9378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9380 = 7'h7a == _myNewVec_56_T_3[6:0] ? myVec_122 : _GEN_9379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9381 = 7'h7b == _myNewVec_56_T_3[6:0] ? myVec_123 : _GEN_9380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9382 = 7'h7c == _myNewVec_56_T_3[6:0] ? myVec_124 : _GEN_9381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9383 = 7'h7d == _myNewVec_56_T_3[6:0] ? myVec_125 : _GEN_9382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9384 = 7'h7e == _myNewVec_56_T_3[6:0] ? myVec_126 : _GEN_9383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_56 = 7'h7f == _myNewVec_56_T_3[6:0] ? myVec_127 : _GEN_9384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_55_T_3 = _myNewVec_127_T_1 + 16'h48; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_9387 = 7'h1 == _myNewVec_55_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9388 = 7'h2 == _myNewVec_55_T_3[6:0] ? myVec_2 : _GEN_9387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9389 = 7'h3 == _myNewVec_55_T_3[6:0] ? myVec_3 : _GEN_9388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9390 = 7'h4 == _myNewVec_55_T_3[6:0] ? myVec_4 : _GEN_9389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9391 = 7'h5 == _myNewVec_55_T_3[6:0] ? myVec_5 : _GEN_9390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9392 = 7'h6 == _myNewVec_55_T_3[6:0] ? myVec_6 : _GEN_9391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9393 = 7'h7 == _myNewVec_55_T_3[6:0] ? myVec_7 : _GEN_9392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9394 = 7'h8 == _myNewVec_55_T_3[6:0] ? myVec_8 : _GEN_9393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9395 = 7'h9 == _myNewVec_55_T_3[6:0] ? myVec_9 : _GEN_9394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9396 = 7'ha == _myNewVec_55_T_3[6:0] ? myVec_10 : _GEN_9395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9397 = 7'hb == _myNewVec_55_T_3[6:0] ? myVec_11 : _GEN_9396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9398 = 7'hc == _myNewVec_55_T_3[6:0] ? myVec_12 : _GEN_9397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9399 = 7'hd == _myNewVec_55_T_3[6:0] ? myVec_13 : _GEN_9398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9400 = 7'he == _myNewVec_55_T_3[6:0] ? myVec_14 : _GEN_9399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9401 = 7'hf == _myNewVec_55_T_3[6:0] ? myVec_15 : _GEN_9400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9402 = 7'h10 == _myNewVec_55_T_3[6:0] ? myVec_16 : _GEN_9401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9403 = 7'h11 == _myNewVec_55_T_3[6:0] ? myVec_17 : _GEN_9402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9404 = 7'h12 == _myNewVec_55_T_3[6:0] ? myVec_18 : _GEN_9403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9405 = 7'h13 == _myNewVec_55_T_3[6:0] ? myVec_19 : _GEN_9404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9406 = 7'h14 == _myNewVec_55_T_3[6:0] ? myVec_20 : _GEN_9405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9407 = 7'h15 == _myNewVec_55_T_3[6:0] ? myVec_21 : _GEN_9406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9408 = 7'h16 == _myNewVec_55_T_3[6:0] ? myVec_22 : _GEN_9407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9409 = 7'h17 == _myNewVec_55_T_3[6:0] ? myVec_23 : _GEN_9408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9410 = 7'h18 == _myNewVec_55_T_3[6:0] ? myVec_24 : _GEN_9409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9411 = 7'h19 == _myNewVec_55_T_3[6:0] ? myVec_25 : _GEN_9410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9412 = 7'h1a == _myNewVec_55_T_3[6:0] ? myVec_26 : _GEN_9411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9413 = 7'h1b == _myNewVec_55_T_3[6:0] ? myVec_27 : _GEN_9412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9414 = 7'h1c == _myNewVec_55_T_3[6:0] ? myVec_28 : _GEN_9413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9415 = 7'h1d == _myNewVec_55_T_3[6:0] ? myVec_29 : _GEN_9414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9416 = 7'h1e == _myNewVec_55_T_3[6:0] ? myVec_30 : _GEN_9415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9417 = 7'h1f == _myNewVec_55_T_3[6:0] ? myVec_31 : _GEN_9416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9418 = 7'h20 == _myNewVec_55_T_3[6:0] ? myVec_32 : _GEN_9417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9419 = 7'h21 == _myNewVec_55_T_3[6:0] ? myVec_33 : _GEN_9418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9420 = 7'h22 == _myNewVec_55_T_3[6:0] ? myVec_34 : _GEN_9419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9421 = 7'h23 == _myNewVec_55_T_3[6:0] ? myVec_35 : _GEN_9420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9422 = 7'h24 == _myNewVec_55_T_3[6:0] ? myVec_36 : _GEN_9421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9423 = 7'h25 == _myNewVec_55_T_3[6:0] ? myVec_37 : _GEN_9422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9424 = 7'h26 == _myNewVec_55_T_3[6:0] ? myVec_38 : _GEN_9423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9425 = 7'h27 == _myNewVec_55_T_3[6:0] ? myVec_39 : _GEN_9424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9426 = 7'h28 == _myNewVec_55_T_3[6:0] ? myVec_40 : _GEN_9425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9427 = 7'h29 == _myNewVec_55_T_3[6:0] ? myVec_41 : _GEN_9426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9428 = 7'h2a == _myNewVec_55_T_3[6:0] ? myVec_42 : _GEN_9427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9429 = 7'h2b == _myNewVec_55_T_3[6:0] ? myVec_43 : _GEN_9428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9430 = 7'h2c == _myNewVec_55_T_3[6:0] ? myVec_44 : _GEN_9429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9431 = 7'h2d == _myNewVec_55_T_3[6:0] ? myVec_45 : _GEN_9430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9432 = 7'h2e == _myNewVec_55_T_3[6:0] ? myVec_46 : _GEN_9431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9433 = 7'h2f == _myNewVec_55_T_3[6:0] ? myVec_47 : _GEN_9432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9434 = 7'h30 == _myNewVec_55_T_3[6:0] ? myVec_48 : _GEN_9433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9435 = 7'h31 == _myNewVec_55_T_3[6:0] ? myVec_49 : _GEN_9434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9436 = 7'h32 == _myNewVec_55_T_3[6:0] ? myVec_50 : _GEN_9435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9437 = 7'h33 == _myNewVec_55_T_3[6:0] ? myVec_51 : _GEN_9436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9438 = 7'h34 == _myNewVec_55_T_3[6:0] ? myVec_52 : _GEN_9437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9439 = 7'h35 == _myNewVec_55_T_3[6:0] ? myVec_53 : _GEN_9438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9440 = 7'h36 == _myNewVec_55_T_3[6:0] ? myVec_54 : _GEN_9439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9441 = 7'h37 == _myNewVec_55_T_3[6:0] ? myVec_55 : _GEN_9440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9442 = 7'h38 == _myNewVec_55_T_3[6:0] ? myVec_56 : _GEN_9441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9443 = 7'h39 == _myNewVec_55_T_3[6:0] ? myVec_57 : _GEN_9442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9444 = 7'h3a == _myNewVec_55_T_3[6:0] ? myVec_58 : _GEN_9443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9445 = 7'h3b == _myNewVec_55_T_3[6:0] ? myVec_59 : _GEN_9444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9446 = 7'h3c == _myNewVec_55_T_3[6:0] ? myVec_60 : _GEN_9445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9447 = 7'h3d == _myNewVec_55_T_3[6:0] ? myVec_61 : _GEN_9446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9448 = 7'h3e == _myNewVec_55_T_3[6:0] ? myVec_62 : _GEN_9447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9449 = 7'h3f == _myNewVec_55_T_3[6:0] ? myVec_63 : _GEN_9448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9450 = 7'h40 == _myNewVec_55_T_3[6:0] ? myVec_64 : _GEN_9449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9451 = 7'h41 == _myNewVec_55_T_3[6:0] ? myVec_65 : _GEN_9450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9452 = 7'h42 == _myNewVec_55_T_3[6:0] ? myVec_66 : _GEN_9451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9453 = 7'h43 == _myNewVec_55_T_3[6:0] ? myVec_67 : _GEN_9452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9454 = 7'h44 == _myNewVec_55_T_3[6:0] ? myVec_68 : _GEN_9453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9455 = 7'h45 == _myNewVec_55_T_3[6:0] ? myVec_69 : _GEN_9454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9456 = 7'h46 == _myNewVec_55_T_3[6:0] ? myVec_70 : _GEN_9455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9457 = 7'h47 == _myNewVec_55_T_3[6:0] ? myVec_71 : _GEN_9456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9458 = 7'h48 == _myNewVec_55_T_3[6:0] ? myVec_72 : _GEN_9457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9459 = 7'h49 == _myNewVec_55_T_3[6:0] ? myVec_73 : _GEN_9458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9460 = 7'h4a == _myNewVec_55_T_3[6:0] ? myVec_74 : _GEN_9459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9461 = 7'h4b == _myNewVec_55_T_3[6:0] ? myVec_75 : _GEN_9460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9462 = 7'h4c == _myNewVec_55_T_3[6:0] ? myVec_76 : _GEN_9461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9463 = 7'h4d == _myNewVec_55_T_3[6:0] ? myVec_77 : _GEN_9462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9464 = 7'h4e == _myNewVec_55_T_3[6:0] ? myVec_78 : _GEN_9463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9465 = 7'h4f == _myNewVec_55_T_3[6:0] ? myVec_79 : _GEN_9464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9466 = 7'h50 == _myNewVec_55_T_3[6:0] ? myVec_80 : _GEN_9465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9467 = 7'h51 == _myNewVec_55_T_3[6:0] ? myVec_81 : _GEN_9466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9468 = 7'h52 == _myNewVec_55_T_3[6:0] ? myVec_82 : _GEN_9467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9469 = 7'h53 == _myNewVec_55_T_3[6:0] ? myVec_83 : _GEN_9468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9470 = 7'h54 == _myNewVec_55_T_3[6:0] ? myVec_84 : _GEN_9469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9471 = 7'h55 == _myNewVec_55_T_3[6:0] ? myVec_85 : _GEN_9470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9472 = 7'h56 == _myNewVec_55_T_3[6:0] ? myVec_86 : _GEN_9471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9473 = 7'h57 == _myNewVec_55_T_3[6:0] ? myVec_87 : _GEN_9472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9474 = 7'h58 == _myNewVec_55_T_3[6:0] ? myVec_88 : _GEN_9473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9475 = 7'h59 == _myNewVec_55_T_3[6:0] ? myVec_89 : _GEN_9474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9476 = 7'h5a == _myNewVec_55_T_3[6:0] ? myVec_90 : _GEN_9475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9477 = 7'h5b == _myNewVec_55_T_3[6:0] ? myVec_91 : _GEN_9476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9478 = 7'h5c == _myNewVec_55_T_3[6:0] ? myVec_92 : _GEN_9477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9479 = 7'h5d == _myNewVec_55_T_3[6:0] ? myVec_93 : _GEN_9478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9480 = 7'h5e == _myNewVec_55_T_3[6:0] ? myVec_94 : _GEN_9479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9481 = 7'h5f == _myNewVec_55_T_3[6:0] ? myVec_95 : _GEN_9480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9482 = 7'h60 == _myNewVec_55_T_3[6:0] ? myVec_96 : _GEN_9481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9483 = 7'h61 == _myNewVec_55_T_3[6:0] ? myVec_97 : _GEN_9482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9484 = 7'h62 == _myNewVec_55_T_3[6:0] ? myVec_98 : _GEN_9483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9485 = 7'h63 == _myNewVec_55_T_3[6:0] ? myVec_99 : _GEN_9484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9486 = 7'h64 == _myNewVec_55_T_3[6:0] ? myVec_100 : _GEN_9485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9487 = 7'h65 == _myNewVec_55_T_3[6:0] ? myVec_101 : _GEN_9486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9488 = 7'h66 == _myNewVec_55_T_3[6:0] ? myVec_102 : _GEN_9487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9489 = 7'h67 == _myNewVec_55_T_3[6:0] ? myVec_103 : _GEN_9488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9490 = 7'h68 == _myNewVec_55_T_3[6:0] ? myVec_104 : _GEN_9489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9491 = 7'h69 == _myNewVec_55_T_3[6:0] ? myVec_105 : _GEN_9490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9492 = 7'h6a == _myNewVec_55_T_3[6:0] ? myVec_106 : _GEN_9491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9493 = 7'h6b == _myNewVec_55_T_3[6:0] ? myVec_107 : _GEN_9492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9494 = 7'h6c == _myNewVec_55_T_3[6:0] ? myVec_108 : _GEN_9493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9495 = 7'h6d == _myNewVec_55_T_3[6:0] ? myVec_109 : _GEN_9494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9496 = 7'h6e == _myNewVec_55_T_3[6:0] ? myVec_110 : _GEN_9495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9497 = 7'h6f == _myNewVec_55_T_3[6:0] ? myVec_111 : _GEN_9496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9498 = 7'h70 == _myNewVec_55_T_3[6:0] ? myVec_112 : _GEN_9497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9499 = 7'h71 == _myNewVec_55_T_3[6:0] ? myVec_113 : _GEN_9498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9500 = 7'h72 == _myNewVec_55_T_3[6:0] ? myVec_114 : _GEN_9499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9501 = 7'h73 == _myNewVec_55_T_3[6:0] ? myVec_115 : _GEN_9500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9502 = 7'h74 == _myNewVec_55_T_3[6:0] ? myVec_116 : _GEN_9501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9503 = 7'h75 == _myNewVec_55_T_3[6:0] ? myVec_117 : _GEN_9502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9504 = 7'h76 == _myNewVec_55_T_3[6:0] ? myVec_118 : _GEN_9503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9505 = 7'h77 == _myNewVec_55_T_3[6:0] ? myVec_119 : _GEN_9504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9506 = 7'h78 == _myNewVec_55_T_3[6:0] ? myVec_120 : _GEN_9505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9507 = 7'h79 == _myNewVec_55_T_3[6:0] ? myVec_121 : _GEN_9506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9508 = 7'h7a == _myNewVec_55_T_3[6:0] ? myVec_122 : _GEN_9507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9509 = 7'h7b == _myNewVec_55_T_3[6:0] ? myVec_123 : _GEN_9508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9510 = 7'h7c == _myNewVec_55_T_3[6:0] ? myVec_124 : _GEN_9509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9511 = 7'h7d == _myNewVec_55_T_3[6:0] ? myVec_125 : _GEN_9510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9512 = 7'h7e == _myNewVec_55_T_3[6:0] ? myVec_126 : _GEN_9511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_55 = 7'h7f == _myNewVec_55_T_3[6:0] ? myVec_127 : _GEN_9512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_54_T_3 = _myNewVec_127_T_1 + 16'h49; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_9515 = 7'h1 == _myNewVec_54_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9516 = 7'h2 == _myNewVec_54_T_3[6:0] ? myVec_2 : _GEN_9515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9517 = 7'h3 == _myNewVec_54_T_3[6:0] ? myVec_3 : _GEN_9516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9518 = 7'h4 == _myNewVec_54_T_3[6:0] ? myVec_4 : _GEN_9517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9519 = 7'h5 == _myNewVec_54_T_3[6:0] ? myVec_5 : _GEN_9518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9520 = 7'h6 == _myNewVec_54_T_3[6:0] ? myVec_6 : _GEN_9519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9521 = 7'h7 == _myNewVec_54_T_3[6:0] ? myVec_7 : _GEN_9520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9522 = 7'h8 == _myNewVec_54_T_3[6:0] ? myVec_8 : _GEN_9521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9523 = 7'h9 == _myNewVec_54_T_3[6:0] ? myVec_9 : _GEN_9522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9524 = 7'ha == _myNewVec_54_T_3[6:0] ? myVec_10 : _GEN_9523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9525 = 7'hb == _myNewVec_54_T_3[6:0] ? myVec_11 : _GEN_9524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9526 = 7'hc == _myNewVec_54_T_3[6:0] ? myVec_12 : _GEN_9525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9527 = 7'hd == _myNewVec_54_T_3[6:0] ? myVec_13 : _GEN_9526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9528 = 7'he == _myNewVec_54_T_3[6:0] ? myVec_14 : _GEN_9527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9529 = 7'hf == _myNewVec_54_T_3[6:0] ? myVec_15 : _GEN_9528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9530 = 7'h10 == _myNewVec_54_T_3[6:0] ? myVec_16 : _GEN_9529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9531 = 7'h11 == _myNewVec_54_T_3[6:0] ? myVec_17 : _GEN_9530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9532 = 7'h12 == _myNewVec_54_T_3[6:0] ? myVec_18 : _GEN_9531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9533 = 7'h13 == _myNewVec_54_T_3[6:0] ? myVec_19 : _GEN_9532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9534 = 7'h14 == _myNewVec_54_T_3[6:0] ? myVec_20 : _GEN_9533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9535 = 7'h15 == _myNewVec_54_T_3[6:0] ? myVec_21 : _GEN_9534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9536 = 7'h16 == _myNewVec_54_T_3[6:0] ? myVec_22 : _GEN_9535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9537 = 7'h17 == _myNewVec_54_T_3[6:0] ? myVec_23 : _GEN_9536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9538 = 7'h18 == _myNewVec_54_T_3[6:0] ? myVec_24 : _GEN_9537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9539 = 7'h19 == _myNewVec_54_T_3[6:0] ? myVec_25 : _GEN_9538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9540 = 7'h1a == _myNewVec_54_T_3[6:0] ? myVec_26 : _GEN_9539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9541 = 7'h1b == _myNewVec_54_T_3[6:0] ? myVec_27 : _GEN_9540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9542 = 7'h1c == _myNewVec_54_T_3[6:0] ? myVec_28 : _GEN_9541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9543 = 7'h1d == _myNewVec_54_T_3[6:0] ? myVec_29 : _GEN_9542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9544 = 7'h1e == _myNewVec_54_T_3[6:0] ? myVec_30 : _GEN_9543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9545 = 7'h1f == _myNewVec_54_T_3[6:0] ? myVec_31 : _GEN_9544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9546 = 7'h20 == _myNewVec_54_T_3[6:0] ? myVec_32 : _GEN_9545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9547 = 7'h21 == _myNewVec_54_T_3[6:0] ? myVec_33 : _GEN_9546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9548 = 7'h22 == _myNewVec_54_T_3[6:0] ? myVec_34 : _GEN_9547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9549 = 7'h23 == _myNewVec_54_T_3[6:0] ? myVec_35 : _GEN_9548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9550 = 7'h24 == _myNewVec_54_T_3[6:0] ? myVec_36 : _GEN_9549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9551 = 7'h25 == _myNewVec_54_T_3[6:0] ? myVec_37 : _GEN_9550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9552 = 7'h26 == _myNewVec_54_T_3[6:0] ? myVec_38 : _GEN_9551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9553 = 7'h27 == _myNewVec_54_T_3[6:0] ? myVec_39 : _GEN_9552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9554 = 7'h28 == _myNewVec_54_T_3[6:0] ? myVec_40 : _GEN_9553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9555 = 7'h29 == _myNewVec_54_T_3[6:0] ? myVec_41 : _GEN_9554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9556 = 7'h2a == _myNewVec_54_T_3[6:0] ? myVec_42 : _GEN_9555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9557 = 7'h2b == _myNewVec_54_T_3[6:0] ? myVec_43 : _GEN_9556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9558 = 7'h2c == _myNewVec_54_T_3[6:0] ? myVec_44 : _GEN_9557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9559 = 7'h2d == _myNewVec_54_T_3[6:0] ? myVec_45 : _GEN_9558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9560 = 7'h2e == _myNewVec_54_T_3[6:0] ? myVec_46 : _GEN_9559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9561 = 7'h2f == _myNewVec_54_T_3[6:0] ? myVec_47 : _GEN_9560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9562 = 7'h30 == _myNewVec_54_T_3[6:0] ? myVec_48 : _GEN_9561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9563 = 7'h31 == _myNewVec_54_T_3[6:0] ? myVec_49 : _GEN_9562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9564 = 7'h32 == _myNewVec_54_T_3[6:0] ? myVec_50 : _GEN_9563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9565 = 7'h33 == _myNewVec_54_T_3[6:0] ? myVec_51 : _GEN_9564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9566 = 7'h34 == _myNewVec_54_T_3[6:0] ? myVec_52 : _GEN_9565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9567 = 7'h35 == _myNewVec_54_T_3[6:0] ? myVec_53 : _GEN_9566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9568 = 7'h36 == _myNewVec_54_T_3[6:0] ? myVec_54 : _GEN_9567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9569 = 7'h37 == _myNewVec_54_T_3[6:0] ? myVec_55 : _GEN_9568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9570 = 7'h38 == _myNewVec_54_T_3[6:0] ? myVec_56 : _GEN_9569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9571 = 7'h39 == _myNewVec_54_T_3[6:0] ? myVec_57 : _GEN_9570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9572 = 7'h3a == _myNewVec_54_T_3[6:0] ? myVec_58 : _GEN_9571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9573 = 7'h3b == _myNewVec_54_T_3[6:0] ? myVec_59 : _GEN_9572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9574 = 7'h3c == _myNewVec_54_T_3[6:0] ? myVec_60 : _GEN_9573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9575 = 7'h3d == _myNewVec_54_T_3[6:0] ? myVec_61 : _GEN_9574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9576 = 7'h3e == _myNewVec_54_T_3[6:0] ? myVec_62 : _GEN_9575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9577 = 7'h3f == _myNewVec_54_T_3[6:0] ? myVec_63 : _GEN_9576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9578 = 7'h40 == _myNewVec_54_T_3[6:0] ? myVec_64 : _GEN_9577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9579 = 7'h41 == _myNewVec_54_T_3[6:0] ? myVec_65 : _GEN_9578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9580 = 7'h42 == _myNewVec_54_T_3[6:0] ? myVec_66 : _GEN_9579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9581 = 7'h43 == _myNewVec_54_T_3[6:0] ? myVec_67 : _GEN_9580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9582 = 7'h44 == _myNewVec_54_T_3[6:0] ? myVec_68 : _GEN_9581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9583 = 7'h45 == _myNewVec_54_T_3[6:0] ? myVec_69 : _GEN_9582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9584 = 7'h46 == _myNewVec_54_T_3[6:0] ? myVec_70 : _GEN_9583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9585 = 7'h47 == _myNewVec_54_T_3[6:0] ? myVec_71 : _GEN_9584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9586 = 7'h48 == _myNewVec_54_T_3[6:0] ? myVec_72 : _GEN_9585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9587 = 7'h49 == _myNewVec_54_T_3[6:0] ? myVec_73 : _GEN_9586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9588 = 7'h4a == _myNewVec_54_T_3[6:0] ? myVec_74 : _GEN_9587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9589 = 7'h4b == _myNewVec_54_T_3[6:0] ? myVec_75 : _GEN_9588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9590 = 7'h4c == _myNewVec_54_T_3[6:0] ? myVec_76 : _GEN_9589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9591 = 7'h4d == _myNewVec_54_T_3[6:0] ? myVec_77 : _GEN_9590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9592 = 7'h4e == _myNewVec_54_T_3[6:0] ? myVec_78 : _GEN_9591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9593 = 7'h4f == _myNewVec_54_T_3[6:0] ? myVec_79 : _GEN_9592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9594 = 7'h50 == _myNewVec_54_T_3[6:0] ? myVec_80 : _GEN_9593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9595 = 7'h51 == _myNewVec_54_T_3[6:0] ? myVec_81 : _GEN_9594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9596 = 7'h52 == _myNewVec_54_T_3[6:0] ? myVec_82 : _GEN_9595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9597 = 7'h53 == _myNewVec_54_T_3[6:0] ? myVec_83 : _GEN_9596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9598 = 7'h54 == _myNewVec_54_T_3[6:0] ? myVec_84 : _GEN_9597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9599 = 7'h55 == _myNewVec_54_T_3[6:0] ? myVec_85 : _GEN_9598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9600 = 7'h56 == _myNewVec_54_T_3[6:0] ? myVec_86 : _GEN_9599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9601 = 7'h57 == _myNewVec_54_T_3[6:0] ? myVec_87 : _GEN_9600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9602 = 7'h58 == _myNewVec_54_T_3[6:0] ? myVec_88 : _GEN_9601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9603 = 7'h59 == _myNewVec_54_T_3[6:0] ? myVec_89 : _GEN_9602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9604 = 7'h5a == _myNewVec_54_T_3[6:0] ? myVec_90 : _GEN_9603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9605 = 7'h5b == _myNewVec_54_T_3[6:0] ? myVec_91 : _GEN_9604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9606 = 7'h5c == _myNewVec_54_T_3[6:0] ? myVec_92 : _GEN_9605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9607 = 7'h5d == _myNewVec_54_T_3[6:0] ? myVec_93 : _GEN_9606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9608 = 7'h5e == _myNewVec_54_T_3[6:0] ? myVec_94 : _GEN_9607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9609 = 7'h5f == _myNewVec_54_T_3[6:0] ? myVec_95 : _GEN_9608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9610 = 7'h60 == _myNewVec_54_T_3[6:0] ? myVec_96 : _GEN_9609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9611 = 7'h61 == _myNewVec_54_T_3[6:0] ? myVec_97 : _GEN_9610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9612 = 7'h62 == _myNewVec_54_T_3[6:0] ? myVec_98 : _GEN_9611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9613 = 7'h63 == _myNewVec_54_T_3[6:0] ? myVec_99 : _GEN_9612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9614 = 7'h64 == _myNewVec_54_T_3[6:0] ? myVec_100 : _GEN_9613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9615 = 7'h65 == _myNewVec_54_T_3[6:0] ? myVec_101 : _GEN_9614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9616 = 7'h66 == _myNewVec_54_T_3[6:0] ? myVec_102 : _GEN_9615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9617 = 7'h67 == _myNewVec_54_T_3[6:0] ? myVec_103 : _GEN_9616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9618 = 7'h68 == _myNewVec_54_T_3[6:0] ? myVec_104 : _GEN_9617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9619 = 7'h69 == _myNewVec_54_T_3[6:0] ? myVec_105 : _GEN_9618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9620 = 7'h6a == _myNewVec_54_T_3[6:0] ? myVec_106 : _GEN_9619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9621 = 7'h6b == _myNewVec_54_T_3[6:0] ? myVec_107 : _GEN_9620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9622 = 7'h6c == _myNewVec_54_T_3[6:0] ? myVec_108 : _GEN_9621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9623 = 7'h6d == _myNewVec_54_T_3[6:0] ? myVec_109 : _GEN_9622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9624 = 7'h6e == _myNewVec_54_T_3[6:0] ? myVec_110 : _GEN_9623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9625 = 7'h6f == _myNewVec_54_T_3[6:0] ? myVec_111 : _GEN_9624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9626 = 7'h70 == _myNewVec_54_T_3[6:0] ? myVec_112 : _GEN_9625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9627 = 7'h71 == _myNewVec_54_T_3[6:0] ? myVec_113 : _GEN_9626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9628 = 7'h72 == _myNewVec_54_T_3[6:0] ? myVec_114 : _GEN_9627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9629 = 7'h73 == _myNewVec_54_T_3[6:0] ? myVec_115 : _GEN_9628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9630 = 7'h74 == _myNewVec_54_T_3[6:0] ? myVec_116 : _GEN_9629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9631 = 7'h75 == _myNewVec_54_T_3[6:0] ? myVec_117 : _GEN_9630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9632 = 7'h76 == _myNewVec_54_T_3[6:0] ? myVec_118 : _GEN_9631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9633 = 7'h77 == _myNewVec_54_T_3[6:0] ? myVec_119 : _GEN_9632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9634 = 7'h78 == _myNewVec_54_T_3[6:0] ? myVec_120 : _GEN_9633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9635 = 7'h79 == _myNewVec_54_T_3[6:0] ? myVec_121 : _GEN_9634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9636 = 7'h7a == _myNewVec_54_T_3[6:0] ? myVec_122 : _GEN_9635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9637 = 7'h7b == _myNewVec_54_T_3[6:0] ? myVec_123 : _GEN_9636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9638 = 7'h7c == _myNewVec_54_T_3[6:0] ? myVec_124 : _GEN_9637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9639 = 7'h7d == _myNewVec_54_T_3[6:0] ? myVec_125 : _GEN_9638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9640 = 7'h7e == _myNewVec_54_T_3[6:0] ? myVec_126 : _GEN_9639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_54 = 7'h7f == _myNewVec_54_T_3[6:0] ? myVec_127 : _GEN_9640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_53_T_3 = _myNewVec_127_T_1 + 16'h4a; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_9643 = 7'h1 == _myNewVec_53_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9644 = 7'h2 == _myNewVec_53_T_3[6:0] ? myVec_2 : _GEN_9643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9645 = 7'h3 == _myNewVec_53_T_3[6:0] ? myVec_3 : _GEN_9644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9646 = 7'h4 == _myNewVec_53_T_3[6:0] ? myVec_4 : _GEN_9645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9647 = 7'h5 == _myNewVec_53_T_3[6:0] ? myVec_5 : _GEN_9646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9648 = 7'h6 == _myNewVec_53_T_3[6:0] ? myVec_6 : _GEN_9647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9649 = 7'h7 == _myNewVec_53_T_3[6:0] ? myVec_7 : _GEN_9648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9650 = 7'h8 == _myNewVec_53_T_3[6:0] ? myVec_8 : _GEN_9649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9651 = 7'h9 == _myNewVec_53_T_3[6:0] ? myVec_9 : _GEN_9650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9652 = 7'ha == _myNewVec_53_T_3[6:0] ? myVec_10 : _GEN_9651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9653 = 7'hb == _myNewVec_53_T_3[6:0] ? myVec_11 : _GEN_9652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9654 = 7'hc == _myNewVec_53_T_3[6:0] ? myVec_12 : _GEN_9653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9655 = 7'hd == _myNewVec_53_T_3[6:0] ? myVec_13 : _GEN_9654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9656 = 7'he == _myNewVec_53_T_3[6:0] ? myVec_14 : _GEN_9655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9657 = 7'hf == _myNewVec_53_T_3[6:0] ? myVec_15 : _GEN_9656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9658 = 7'h10 == _myNewVec_53_T_3[6:0] ? myVec_16 : _GEN_9657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9659 = 7'h11 == _myNewVec_53_T_3[6:0] ? myVec_17 : _GEN_9658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9660 = 7'h12 == _myNewVec_53_T_3[6:0] ? myVec_18 : _GEN_9659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9661 = 7'h13 == _myNewVec_53_T_3[6:0] ? myVec_19 : _GEN_9660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9662 = 7'h14 == _myNewVec_53_T_3[6:0] ? myVec_20 : _GEN_9661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9663 = 7'h15 == _myNewVec_53_T_3[6:0] ? myVec_21 : _GEN_9662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9664 = 7'h16 == _myNewVec_53_T_3[6:0] ? myVec_22 : _GEN_9663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9665 = 7'h17 == _myNewVec_53_T_3[6:0] ? myVec_23 : _GEN_9664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9666 = 7'h18 == _myNewVec_53_T_3[6:0] ? myVec_24 : _GEN_9665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9667 = 7'h19 == _myNewVec_53_T_3[6:0] ? myVec_25 : _GEN_9666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9668 = 7'h1a == _myNewVec_53_T_3[6:0] ? myVec_26 : _GEN_9667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9669 = 7'h1b == _myNewVec_53_T_3[6:0] ? myVec_27 : _GEN_9668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9670 = 7'h1c == _myNewVec_53_T_3[6:0] ? myVec_28 : _GEN_9669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9671 = 7'h1d == _myNewVec_53_T_3[6:0] ? myVec_29 : _GEN_9670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9672 = 7'h1e == _myNewVec_53_T_3[6:0] ? myVec_30 : _GEN_9671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9673 = 7'h1f == _myNewVec_53_T_3[6:0] ? myVec_31 : _GEN_9672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9674 = 7'h20 == _myNewVec_53_T_3[6:0] ? myVec_32 : _GEN_9673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9675 = 7'h21 == _myNewVec_53_T_3[6:0] ? myVec_33 : _GEN_9674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9676 = 7'h22 == _myNewVec_53_T_3[6:0] ? myVec_34 : _GEN_9675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9677 = 7'h23 == _myNewVec_53_T_3[6:0] ? myVec_35 : _GEN_9676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9678 = 7'h24 == _myNewVec_53_T_3[6:0] ? myVec_36 : _GEN_9677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9679 = 7'h25 == _myNewVec_53_T_3[6:0] ? myVec_37 : _GEN_9678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9680 = 7'h26 == _myNewVec_53_T_3[6:0] ? myVec_38 : _GEN_9679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9681 = 7'h27 == _myNewVec_53_T_3[6:0] ? myVec_39 : _GEN_9680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9682 = 7'h28 == _myNewVec_53_T_3[6:0] ? myVec_40 : _GEN_9681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9683 = 7'h29 == _myNewVec_53_T_3[6:0] ? myVec_41 : _GEN_9682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9684 = 7'h2a == _myNewVec_53_T_3[6:0] ? myVec_42 : _GEN_9683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9685 = 7'h2b == _myNewVec_53_T_3[6:0] ? myVec_43 : _GEN_9684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9686 = 7'h2c == _myNewVec_53_T_3[6:0] ? myVec_44 : _GEN_9685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9687 = 7'h2d == _myNewVec_53_T_3[6:0] ? myVec_45 : _GEN_9686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9688 = 7'h2e == _myNewVec_53_T_3[6:0] ? myVec_46 : _GEN_9687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9689 = 7'h2f == _myNewVec_53_T_3[6:0] ? myVec_47 : _GEN_9688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9690 = 7'h30 == _myNewVec_53_T_3[6:0] ? myVec_48 : _GEN_9689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9691 = 7'h31 == _myNewVec_53_T_3[6:0] ? myVec_49 : _GEN_9690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9692 = 7'h32 == _myNewVec_53_T_3[6:0] ? myVec_50 : _GEN_9691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9693 = 7'h33 == _myNewVec_53_T_3[6:0] ? myVec_51 : _GEN_9692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9694 = 7'h34 == _myNewVec_53_T_3[6:0] ? myVec_52 : _GEN_9693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9695 = 7'h35 == _myNewVec_53_T_3[6:0] ? myVec_53 : _GEN_9694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9696 = 7'h36 == _myNewVec_53_T_3[6:0] ? myVec_54 : _GEN_9695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9697 = 7'h37 == _myNewVec_53_T_3[6:0] ? myVec_55 : _GEN_9696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9698 = 7'h38 == _myNewVec_53_T_3[6:0] ? myVec_56 : _GEN_9697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9699 = 7'h39 == _myNewVec_53_T_3[6:0] ? myVec_57 : _GEN_9698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9700 = 7'h3a == _myNewVec_53_T_3[6:0] ? myVec_58 : _GEN_9699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9701 = 7'h3b == _myNewVec_53_T_3[6:0] ? myVec_59 : _GEN_9700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9702 = 7'h3c == _myNewVec_53_T_3[6:0] ? myVec_60 : _GEN_9701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9703 = 7'h3d == _myNewVec_53_T_3[6:0] ? myVec_61 : _GEN_9702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9704 = 7'h3e == _myNewVec_53_T_3[6:0] ? myVec_62 : _GEN_9703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9705 = 7'h3f == _myNewVec_53_T_3[6:0] ? myVec_63 : _GEN_9704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9706 = 7'h40 == _myNewVec_53_T_3[6:0] ? myVec_64 : _GEN_9705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9707 = 7'h41 == _myNewVec_53_T_3[6:0] ? myVec_65 : _GEN_9706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9708 = 7'h42 == _myNewVec_53_T_3[6:0] ? myVec_66 : _GEN_9707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9709 = 7'h43 == _myNewVec_53_T_3[6:0] ? myVec_67 : _GEN_9708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9710 = 7'h44 == _myNewVec_53_T_3[6:0] ? myVec_68 : _GEN_9709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9711 = 7'h45 == _myNewVec_53_T_3[6:0] ? myVec_69 : _GEN_9710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9712 = 7'h46 == _myNewVec_53_T_3[6:0] ? myVec_70 : _GEN_9711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9713 = 7'h47 == _myNewVec_53_T_3[6:0] ? myVec_71 : _GEN_9712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9714 = 7'h48 == _myNewVec_53_T_3[6:0] ? myVec_72 : _GEN_9713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9715 = 7'h49 == _myNewVec_53_T_3[6:0] ? myVec_73 : _GEN_9714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9716 = 7'h4a == _myNewVec_53_T_3[6:0] ? myVec_74 : _GEN_9715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9717 = 7'h4b == _myNewVec_53_T_3[6:0] ? myVec_75 : _GEN_9716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9718 = 7'h4c == _myNewVec_53_T_3[6:0] ? myVec_76 : _GEN_9717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9719 = 7'h4d == _myNewVec_53_T_3[6:0] ? myVec_77 : _GEN_9718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9720 = 7'h4e == _myNewVec_53_T_3[6:0] ? myVec_78 : _GEN_9719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9721 = 7'h4f == _myNewVec_53_T_3[6:0] ? myVec_79 : _GEN_9720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9722 = 7'h50 == _myNewVec_53_T_3[6:0] ? myVec_80 : _GEN_9721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9723 = 7'h51 == _myNewVec_53_T_3[6:0] ? myVec_81 : _GEN_9722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9724 = 7'h52 == _myNewVec_53_T_3[6:0] ? myVec_82 : _GEN_9723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9725 = 7'h53 == _myNewVec_53_T_3[6:0] ? myVec_83 : _GEN_9724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9726 = 7'h54 == _myNewVec_53_T_3[6:0] ? myVec_84 : _GEN_9725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9727 = 7'h55 == _myNewVec_53_T_3[6:0] ? myVec_85 : _GEN_9726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9728 = 7'h56 == _myNewVec_53_T_3[6:0] ? myVec_86 : _GEN_9727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9729 = 7'h57 == _myNewVec_53_T_3[6:0] ? myVec_87 : _GEN_9728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9730 = 7'h58 == _myNewVec_53_T_3[6:0] ? myVec_88 : _GEN_9729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9731 = 7'h59 == _myNewVec_53_T_3[6:0] ? myVec_89 : _GEN_9730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9732 = 7'h5a == _myNewVec_53_T_3[6:0] ? myVec_90 : _GEN_9731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9733 = 7'h5b == _myNewVec_53_T_3[6:0] ? myVec_91 : _GEN_9732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9734 = 7'h5c == _myNewVec_53_T_3[6:0] ? myVec_92 : _GEN_9733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9735 = 7'h5d == _myNewVec_53_T_3[6:0] ? myVec_93 : _GEN_9734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9736 = 7'h5e == _myNewVec_53_T_3[6:0] ? myVec_94 : _GEN_9735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9737 = 7'h5f == _myNewVec_53_T_3[6:0] ? myVec_95 : _GEN_9736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9738 = 7'h60 == _myNewVec_53_T_3[6:0] ? myVec_96 : _GEN_9737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9739 = 7'h61 == _myNewVec_53_T_3[6:0] ? myVec_97 : _GEN_9738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9740 = 7'h62 == _myNewVec_53_T_3[6:0] ? myVec_98 : _GEN_9739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9741 = 7'h63 == _myNewVec_53_T_3[6:0] ? myVec_99 : _GEN_9740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9742 = 7'h64 == _myNewVec_53_T_3[6:0] ? myVec_100 : _GEN_9741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9743 = 7'h65 == _myNewVec_53_T_3[6:0] ? myVec_101 : _GEN_9742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9744 = 7'h66 == _myNewVec_53_T_3[6:0] ? myVec_102 : _GEN_9743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9745 = 7'h67 == _myNewVec_53_T_3[6:0] ? myVec_103 : _GEN_9744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9746 = 7'h68 == _myNewVec_53_T_3[6:0] ? myVec_104 : _GEN_9745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9747 = 7'h69 == _myNewVec_53_T_3[6:0] ? myVec_105 : _GEN_9746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9748 = 7'h6a == _myNewVec_53_T_3[6:0] ? myVec_106 : _GEN_9747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9749 = 7'h6b == _myNewVec_53_T_3[6:0] ? myVec_107 : _GEN_9748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9750 = 7'h6c == _myNewVec_53_T_3[6:0] ? myVec_108 : _GEN_9749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9751 = 7'h6d == _myNewVec_53_T_3[6:0] ? myVec_109 : _GEN_9750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9752 = 7'h6e == _myNewVec_53_T_3[6:0] ? myVec_110 : _GEN_9751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9753 = 7'h6f == _myNewVec_53_T_3[6:0] ? myVec_111 : _GEN_9752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9754 = 7'h70 == _myNewVec_53_T_3[6:0] ? myVec_112 : _GEN_9753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9755 = 7'h71 == _myNewVec_53_T_3[6:0] ? myVec_113 : _GEN_9754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9756 = 7'h72 == _myNewVec_53_T_3[6:0] ? myVec_114 : _GEN_9755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9757 = 7'h73 == _myNewVec_53_T_3[6:0] ? myVec_115 : _GEN_9756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9758 = 7'h74 == _myNewVec_53_T_3[6:0] ? myVec_116 : _GEN_9757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9759 = 7'h75 == _myNewVec_53_T_3[6:0] ? myVec_117 : _GEN_9758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9760 = 7'h76 == _myNewVec_53_T_3[6:0] ? myVec_118 : _GEN_9759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9761 = 7'h77 == _myNewVec_53_T_3[6:0] ? myVec_119 : _GEN_9760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9762 = 7'h78 == _myNewVec_53_T_3[6:0] ? myVec_120 : _GEN_9761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9763 = 7'h79 == _myNewVec_53_T_3[6:0] ? myVec_121 : _GEN_9762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9764 = 7'h7a == _myNewVec_53_T_3[6:0] ? myVec_122 : _GEN_9763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9765 = 7'h7b == _myNewVec_53_T_3[6:0] ? myVec_123 : _GEN_9764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9766 = 7'h7c == _myNewVec_53_T_3[6:0] ? myVec_124 : _GEN_9765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9767 = 7'h7d == _myNewVec_53_T_3[6:0] ? myVec_125 : _GEN_9766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9768 = 7'h7e == _myNewVec_53_T_3[6:0] ? myVec_126 : _GEN_9767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_53 = 7'h7f == _myNewVec_53_T_3[6:0] ? myVec_127 : _GEN_9768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_52_T_3 = _myNewVec_127_T_1 + 16'h4b; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_9771 = 7'h1 == _myNewVec_52_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9772 = 7'h2 == _myNewVec_52_T_3[6:0] ? myVec_2 : _GEN_9771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9773 = 7'h3 == _myNewVec_52_T_3[6:0] ? myVec_3 : _GEN_9772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9774 = 7'h4 == _myNewVec_52_T_3[6:0] ? myVec_4 : _GEN_9773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9775 = 7'h5 == _myNewVec_52_T_3[6:0] ? myVec_5 : _GEN_9774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9776 = 7'h6 == _myNewVec_52_T_3[6:0] ? myVec_6 : _GEN_9775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9777 = 7'h7 == _myNewVec_52_T_3[6:0] ? myVec_7 : _GEN_9776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9778 = 7'h8 == _myNewVec_52_T_3[6:0] ? myVec_8 : _GEN_9777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9779 = 7'h9 == _myNewVec_52_T_3[6:0] ? myVec_9 : _GEN_9778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9780 = 7'ha == _myNewVec_52_T_3[6:0] ? myVec_10 : _GEN_9779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9781 = 7'hb == _myNewVec_52_T_3[6:0] ? myVec_11 : _GEN_9780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9782 = 7'hc == _myNewVec_52_T_3[6:0] ? myVec_12 : _GEN_9781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9783 = 7'hd == _myNewVec_52_T_3[6:0] ? myVec_13 : _GEN_9782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9784 = 7'he == _myNewVec_52_T_3[6:0] ? myVec_14 : _GEN_9783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9785 = 7'hf == _myNewVec_52_T_3[6:0] ? myVec_15 : _GEN_9784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9786 = 7'h10 == _myNewVec_52_T_3[6:0] ? myVec_16 : _GEN_9785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9787 = 7'h11 == _myNewVec_52_T_3[6:0] ? myVec_17 : _GEN_9786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9788 = 7'h12 == _myNewVec_52_T_3[6:0] ? myVec_18 : _GEN_9787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9789 = 7'h13 == _myNewVec_52_T_3[6:0] ? myVec_19 : _GEN_9788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9790 = 7'h14 == _myNewVec_52_T_3[6:0] ? myVec_20 : _GEN_9789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9791 = 7'h15 == _myNewVec_52_T_3[6:0] ? myVec_21 : _GEN_9790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9792 = 7'h16 == _myNewVec_52_T_3[6:0] ? myVec_22 : _GEN_9791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9793 = 7'h17 == _myNewVec_52_T_3[6:0] ? myVec_23 : _GEN_9792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9794 = 7'h18 == _myNewVec_52_T_3[6:0] ? myVec_24 : _GEN_9793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9795 = 7'h19 == _myNewVec_52_T_3[6:0] ? myVec_25 : _GEN_9794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9796 = 7'h1a == _myNewVec_52_T_3[6:0] ? myVec_26 : _GEN_9795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9797 = 7'h1b == _myNewVec_52_T_3[6:0] ? myVec_27 : _GEN_9796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9798 = 7'h1c == _myNewVec_52_T_3[6:0] ? myVec_28 : _GEN_9797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9799 = 7'h1d == _myNewVec_52_T_3[6:0] ? myVec_29 : _GEN_9798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9800 = 7'h1e == _myNewVec_52_T_3[6:0] ? myVec_30 : _GEN_9799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9801 = 7'h1f == _myNewVec_52_T_3[6:0] ? myVec_31 : _GEN_9800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9802 = 7'h20 == _myNewVec_52_T_3[6:0] ? myVec_32 : _GEN_9801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9803 = 7'h21 == _myNewVec_52_T_3[6:0] ? myVec_33 : _GEN_9802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9804 = 7'h22 == _myNewVec_52_T_3[6:0] ? myVec_34 : _GEN_9803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9805 = 7'h23 == _myNewVec_52_T_3[6:0] ? myVec_35 : _GEN_9804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9806 = 7'h24 == _myNewVec_52_T_3[6:0] ? myVec_36 : _GEN_9805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9807 = 7'h25 == _myNewVec_52_T_3[6:0] ? myVec_37 : _GEN_9806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9808 = 7'h26 == _myNewVec_52_T_3[6:0] ? myVec_38 : _GEN_9807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9809 = 7'h27 == _myNewVec_52_T_3[6:0] ? myVec_39 : _GEN_9808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9810 = 7'h28 == _myNewVec_52_T_3[6:0] ? myVec_40 : _GEN_9809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9811 = 7'h29 == _myNewVec_52_T_3[6:0] ? myVec_41 : _GEN_9810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9812 = 7'h2a == _myNewVec_52_T_3[6:0] ? myVec_42 : _GEN_9811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9813 = 7'h2b == _myNewVec_52_T_3[6:0] ? myVec_43 : _GEN_9812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9814 = 7'h2c == _myNewVec_52_T_3[6:0] ? myVec_44 : _GEN_9813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9815 = 7'h2d == _myNewVec_52_T_3[6:0] ? myVec_45 : _GEN_9814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9816 = 7'h2e == _myNewVec_52_T_3[6:0] ? myVec_46 : _GEN_9815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9817 = 7'h2f == _myNewVec_52_T_3[6:0] ? myVec_47 : _GEN_9816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9818 = 7'h30 == _myNewVec_52_T_3[6:0] ? myVec_48 : _GEN_9817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9819 = 7'h31 == _myNewVec_52_T_3[6:0] ? myVec_49 : _GEN_9818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9820 = 7'h32 == _myNewVec_52_T_3[6:0] ? myVec_50 : _GEN_9819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9821 = 7'h33 == _myNewVec_52_T_3[6:0] ? myVec_51 : _GEN_9820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9822 = 7'h34 == _myNewVec_52_T_3[6:0] ? myVec_52 : _GEN_9821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9823 = 7'h35 == _myNewVec_52_T_3[6:0] ? myVec_53 : _GEN_9822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9824 = 7'h36 == _myNewVec_52_T_3[6:0] ? myVec_54 : _GEN_9823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9825 = 7'h37 == _myNewVec_52_T_3[6:0] ? myVec_55 : _GEN_9824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9826 = 7'h38 == _myNewVec_52_T_3[6:0] ? myVec_56 : _GEN_9825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9827 = 7'h39 == _myNewVec_52_T_3[6:0] ? myVec_57 : _GEN_9826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9828 = 7'h3a == _myNewVec_52_T_3[6:0] ? myVec_58 : _GEN_9827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9829 = 7'h3b == _myNewVec_52_T_3[6:0] ? myVec_59 : _GEN_9828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9830 = 7'h3c == _myNewVec_52_T_3[6:0] ? myVec_60 : _GEN_9829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9831 = 7'h3d == _myNewVec_52_T_3[6:0] ? myVec_61 : _GEN_9830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9832 = 7'h3e == _myNewVec_52_T_3[6:0] ? myVec_62 : _GEN_9831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9833 = 7'h3f == _myNewVec_52_T_3[6:0] ? myVec_63 : _GEN_9832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9834 = 7'h40 == _myNewVec_52_T_3[6:0] ? myVec_64 : _GEN_9833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9835 = 7'h41 == _myNewVec_52_T_3[6:0] ? myVec_65 : _GEN_9834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9836 = 7'h42 == _myNewVec_52_T_3[6:0] ? myVec_66 : _GEN_9835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9837 = 7'h43 == _myNewVec_52_T_3[6:0] ? myVec_67 : _GEN_9836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9838 = 7'h44 == _myNewVec_52_T_3[6:0] ? myVec_68 : _GEN_9837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9839 = 7'h45 == _myNewVec_52_T_3[6:0] ? myVec_69 : _GEN_9838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9840 = 7'h46 == _myNewVec_52_T_3[6:0] ? myVec_70 : _GEN_9839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9841 = 7'h47 == _myNewVec_52_T_3[6:0] ? myVec_71 : _GEN_9840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9842 = 7'h48 == _myNewVec_52_T_3[6:0] ? myVec_72 : _GEN_9841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9843 = 7'h49 == _myNewVec_52_T_3[6:0] ? myVec_73 : _GEN_9842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9844 = 7'h4a == _myNewVec_52_T_3[6:0] ? myVec_74 : _GEN_9843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9845 = 7'h4b == _myNewVec_52_T_3[6:0] ? myVec_75 : _GEN_9844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9846 = 7'h4c == _myNewVec_52_T_3[6:0] ? myVec_76 : _GEN_9845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9847 = 7'h4d == _myNewVec_52_T_3[6:0] ? myVec_77 : _GEN_9846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9848 = 7'h4e == _myNewVec_52_T_3[6:0] ? myVec_78 : _GEN_9847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9849 = 7'h4f == _myNewVec_52_T_3[6:0] ? myVec_79 : _GEN_9848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9850 = 7'h50 == _myNewVec_52_T_3[6:0] ? myVec_80 : _GEN_9849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9851 = 7'h51 == _myNewVec_52_T_3[6:0] ? myVec_81 : _GEN_9850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9852 = 7'h52 == _myNewVec_52_T_3[6:0] ? myVec_82 : _GEN_9851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9853 = 7'h53 == _myNewVec_52_T_3[6:0] ? myVec_83 : _GEN_9852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9854 = 7'h54 == _myNewVec_52_T_3[6:0] ? myVec_84 : _GEN_9853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9855 = 7'h55 == _myNewVec_52_T_3[6:0] ? myVec_85 : _GEN_9854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9856 = 7'h56 == _myNewVec_52_T_3[6:0] ? myVec_86 : _GEN_9855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9857 = 7'h57 == _myNewVec_52_T_3[6:0] ? myVec_87 : _GEN_9856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9858 = 7'h58 == _myNewVec_52_T_3[6:0] ? myVec_88 : _GEN_9857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9859 = 7'h59 == _myNewVec_52_T_3[6:0] ? myVec_89 : _GEN_9858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9860 = 7'h5a == _myNewVec_52_T_3[6:0] ? myVec_90 : _GEN_9859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9861 = 7'h5b == _myNewVec_52_T_3[6:0] ? myVec_91 : _GEN_9860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9862 = 7'h5c == _myNewVec_52_T_3[6:0] ? myVec_92 : _GEN_9861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9863 = 7'h5d == _myNewVec_52_T_3[6:0] ? myVec_93 : _GEN_9862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9864 = 7'h5e == _myNewVec_52_T_3[6:0] ? myVec_94 : _GEN_9863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9865 = 7'h5f == _myNewVec_52_T_3[6:0] ? myVec_95 : _GEN_9864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9866 = 7'h60 == _myNewVec_52_T_3[6:0] ? myVec_96 : _GEN_9865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9867 = 7'h61 == _myNewVec_52_T_3[6:0] ? myVec_97 : _GEN_9866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9868 = 7'h62 == _myNewVec_52_T_3[6:0] ? myVec_98 : _GEN_9867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9869 = 7'h63 == _myNewVec_52_T_3[6:0] ? myVec_99 : _GEN_9868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9870 = 7'h64 == _myNewVec_52_T_3[6:0] ? myVec_100 : _GEN_9869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9871 = 7'h65 == _myNewVec_52_T_3[6:0] ? myVec_101 : _GEN_9870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9872 = 7'h66 == _myNewVec_52_T_3[6:0] ? myVec_102 : _GEN_9871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9873 = 7'h67 == _myNewVec_52_T_3[6:0] ? myVec_103 : _GEN_9872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9874 = 7'h68 == _myNewVec_52_T_3[6:0] ? myVec_104 : _GEN_9873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9875 = 7'h69 == _myNewVec_52_T_3[6:0] ? myVec_105 : _GEN_9874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9876 = 7'h6a == _myNewVec_52_T_3[6:0] ? myVec_106 : _GEN_9875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9877 = 7'h6b == _myNewVec_52_T_3[6:0] ? myVec_107 : _GEN_9876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9878 = 7'h6c == _myNewVec_52_T_3[6:0] ? myVec_108 : _GEN_9877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9879 = 7'h6d == _myNewVec_52_T_3[6:0] ? myVec_109 : _GEN_9878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9880 = 7'h6e == _myNewVec_52_T_3[6:0] ? myVec_110 : _GEN_9879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9881 = 7'h6f == _myNewVec_52_T_3[6:0] ? myVec_111 : _GEN_9880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9882 = 7'h70 == _myNewVec_52_T_3[6:0] ? myVec_112 : _GEN_9881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9883 = 7'h71 == _myNewVec_52_T_3[6:0] ? myVec_113 : _GEN_9882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9884 = 7'h72 == _myNewVec_52_T_3[6:0] ? myVec_114 : _GEN_9883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9885 = 7'h73 == _myNewVec_52_T_3[6:0] ? myVec_115 : _GEN_9884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9886 = 7'h74 == _myNewVec_52_T_3[6:0] ? myVec_116 : _GEN_9885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9887 = 7'h75 == _myNewVec_52_T_3[6:0] ? myVec_117 : _GEN_9886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9888 = 7'h76 == _myNewVec_52_T_3[6:0] ? myVec_118 : _GEN_9887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9889 = 7'h77 == _myNewVec_52_T_3[6:0] ? myVec_119 : _GEN_9888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9890 = 7'h78 == _myNewVec_52_T_3[6:0] ? myVec_120 : _GEN_9889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9891 = 7'h79 == _myNewVec_52_T_3[6:0] ? myVec_121 : _GEN_9890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9892 = 7'h7a == _myNewVec_52_T_3[6:0] ? myVec_122 : _GEN_9891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9893 = 7'h7b == _myNewVec_52_T_3[6:0] ? myVec_123 : _GEN_9892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9894 = 7'h7c == _myNewVec_52_T_3[6:0] ? myVec_124 : _GEN_9893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9895 = 7'h7d == _myNewVec_52_T_3[6:0] ? myVec_125 : _GEN_9894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9896 = 7'h7e == _myNewVec_52_T_3[6:0] ? myVec_126 : _GEN_9895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_52 = 7'h7f == _myNewVec_52_T_3[6:0] ? myVec_127 : _GEN_9896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_51_T_3 = _myNewVec_127_T_1 + 16'h4c; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_9899 = 7'h1 == _myNewVec_51_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9900 = 7'h2 == _myNewVec_51_T_3[6:0] ? myVec_2 : _GEN_9899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9901 = 7'h3 == _myNewVec_51_T_3[6:0] ? myVec_3 : _GEN_9900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9902 = 7'h4 == _myNewVec_51_T_3[6:0] ? myVec_4 : _GEN_9901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9903 = 7'h5 == _myNewVec_51_T_3[6:0] ? myVec_5 : _GEN_9902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9904 = 7'h6 == _myNewVec_51_T_3[6:0] ? myVec_6 : _GEN_9903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9905 = 7'h7 == _myNewVec_51_T_3[6:0] ? myVec_7 : _GEN_9904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9906 = 7'h8 == _myNewVec_51_T_3[6:0] ? myVec_8 : _GEN_9905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9907 = 7'h9 == _myNewVec_51_T_3[6:0] ? myVec_9 : _GEN_9906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9908 = 7'ha == _myNewVec_51_T_3[6:0] ? myVec_10 : _GEN_9907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9909 = 7'hb == _myNewVec_51_T_3[6:0] ? myVec_11 : _GEN_9908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9910 = 7'hc == _myNewVec_51_T_3[6:0] ? myVec_12 : _GEN_9909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9911 = 7'hd == _myNewVec_51_T_3[6:0] ? myVec_13 : _GEN_9910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9912 = 7'he == _myNewVec_51_T_3[6:0] ? myVec_14 : _GEN_9911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9913 = 7'hf == _myNewVec_51_T_3[6:0] ? myVec_15 : _GEN_9912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9914 = 7'h10 == _myNewVec_51_T_3[6:0] ? myVec_16 : _GEN_9913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9915 = 7'h11 == _myNewVec_51_T_3[6:0] ? myVec_17 : _GEN_9914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9916 = 7'h12 == _myNewVec_51_T_3[6:0] ? myVec_18 : _GEN_9915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9917 = 7'h13 == _myNewVec_51_T_3[6:0] ? myVec_19 : _GEN_9916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9918 = 7'h14 == _myNewVec_51_T_3[6:0] ? myVec_20 : _GEN_9917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9919 = 7'h15 == _myNewVec_51_T_3[6:0] ? myVec_21 : _GEN_9918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9920 = 7'h16 == _myNewVec_51_T_3[6:0] ? myVec_22 : _GEN_9919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9921 = 7'h17 == _myNewVec_51_T_3[6:0] ? myVec_23 : _GEN_9920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9922 = 7'h18 == _myNewVec_51_T_3[6:0] ? myVec_24 : _GEN_9921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9923 = 7'h19 == _myNewVec_51_T_3[6:0] ? myVec_25 : _GEN_9922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9924 = 7'h1a == _myNewVec_51_T_3[6:0] ? myVec_26 : _GEN_9923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9925 = 7'h1b == _myNewVec_51_T_3[6:0] ? myVec_27 : _GEN_9924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9926 = 7'h1c == _myNewVec_51_T_3[6:0] ? myVec_28 : _GEN_9925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9927 = 7'h1d == _myNewVec_51_T_3[6:0] ? myVec_29 : _GEN_9926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9928 = 7'h1e == _myNewVec_51_T_3[6:0] ? myVec_30 : _GEN_9927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9929 = 7'h1f == _myNewVec_51_T_3[6:0] ? myVec_31 : _GEN_9928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9930 = 7'h20 == _myNewVec_51_T_3[6:0] ? myVec_32 : _GEN_9929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9931 = 7'h21 == _myNewVec_51_T_3[6:0] ? myVec_33 : _GEN_9930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9932 = 7'h22 == _myNewVec_51_T_3[6:0] ? myVec_34 : _GEN_9931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9933 = 7'h23 == _myNewVec_51_T_3[6:0] ? myVec_35 : _GEN_9932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9934 = 7'h24 == _myNewVec_51_T_3[6:0] ? myVec_36 : _GEN_9933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9935 = 7'h25 == _myNewVec_51_T_3[6:0] ? myVec_37 : _GEN_9934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9936 = 7'h26 == _myNewVec_51_T_3[6:0] ? myVec_38 : _GEN_9935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9937 = 7'h27 == _myNewVec_51_T_3[6:0] ? myVec_39 : _GEN_9936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9938 = 7'h28 == _myNewVec_51_T_3[6:0] ? myVec_40 : _GEN_9937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9939 = 7'h29 == _myNewVec_51_T_3[6:0] ? myVec_41 : _GEN_9938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9940 = 7'h2a == _myNewVec_51_T_3[6:0] ? myVec_42 : _GEN_9939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9941 = 7'h2b == _myNewVec_51_T_3[6:0] ? myVec_43 : _GEN_9940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9942 = 7'h2c == _myNewVec_51_T_3[6:0] ? myVec_44 : _GEN_9941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9943 = 7'h2d == _myNewVec_51_T_3[6:0] ? myVec_45 : _GEN_9942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9944 = 7'h2e == _myNewVec_51_T_3[6:0] ? myVec_46 : _GEN_9943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9945 = 7'h2f == _myNewVec_51_T_3[6:0] ? myVec_47 : _GEN_9944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9946 = 7'h30 == _myNewVec_51_T_3[6:0] ? myVec_48 : _GEN_9945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9947 = 7'h31 == _myNewVec_51_T_3[6:0] ? myVec_49 : _GEN_9946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9948 = 7'h32 == _myNewVec_51_T_3[6:0] ? myVec_50 : _GEN_9947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9949 = 7'h33 == _myNewVec_51_T_3[6:0] ? myVec_51 : _GEN_9948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9950 = 7'h34 == _myNewVec_51_T_3[6:0] ? myVec_52 : _GEN_9949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9951 = 7'h35 == _myNewVec_51_T_3[6:0] ? myVec_53 : _GEN_9950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9952 = 7'h36 == _myNewVec_51_T_3[6:0] ? myVec_54 : _GEN_9951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9953 = 7'h37 == _myNewVec_51_T_3[6:0] ? myVec_55 : _GEN_9952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9954 = 7'h38 == _myNewVec_51_T_3[6:0] ? myVec_56 : _GEN_9953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9955 = 7'h39 == _myNewVec_51_T_3[6:0] ? myVec_57 : _GEN_9954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9956 = 7'h3a == _myNewVec_51_T_3[6:0] ? myVec_58 : _GEN_9955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9957 = 7'h3b == _myNewVec_51_T_3[6:0] ? myVec_59 : _GEN_9956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9958 = 7'h3c == _myNewVec_51_T_3[6:0] ? myVec_60 : _GEN_9957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9959 = 7'h3d == _myNewVec_51_T_3[6:0] ? myVec_61 : _GEN_9958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9960 = 7'h3e == _myNewVec_51_T_3[6:0] ? myVec_62 : _GEN_9959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9961 = 7'h3f == _myNewVec_51_T_3[6:0] ? myVec_63 : _GEN_9960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9962 = 7'h40 == _myNewVec_51_T_3[6:0] ? myVec_64 : _GEN_9961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9963 = 7'h41 == _myNewVec_51_T_3[6:0] ? myVec_65 : _GEN_9962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9964 = 7'h42 == _myNewVec_51_T_3[6:0] ? myVec_66 : _GEN_9963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9965 = 7'h43 == _myNewVec_51_T_3[6:0] ? myVec_67 : _GEN_9964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9966 = 7'h44 == _myNewVec_51_T_3[6:0] ? myVec_68 : _GEN_9965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9967 = 7'h45 == _myNewVec_51_T_3[6:0] ? myVec_69 : _GEN_9966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9968 = 7'h46 == _myNewVec_51_T_3[6:0] ? myVec_70 : _GEN_9967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9969 = 7'h47 == _myNewVec_51_T_3[6:0] ? myVec_71 : _GEN_9968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9970 = 7'h48 == _myNewVec_51_T_3[6:0] ? myVec_72 : _GEN_9969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9971 = 7'h49 == _myNewVec_51_T_3[6:0] ? myVec_73 : _GEN_9970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9972 = 7'h4a == _myNewVec_51_T_3[6:0] ? myVec_74 : _GEN_9971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9973 = 7'h4b == _myNewVec_51_T_3[6:0] ? myVec_75 : _GEN_9972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9974 = 7'h4c == _myNewVec_51_T_3[6:0] ? myVec_76 : _GEN_9973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9975 = 7'h4d == _myNewVec_51_T_3[6:0] ? myVec_77 : _GEN_9974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9976 = 7'h4e == _myNewVec_51_T_3[6:0] ? myVec_78 : _GEN_9975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9977 = 7'h4f == _myNewVec_51_T_3[6:0] ? myVec_79 : _GEN_9976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9978 = 7'h50 == _myNewVec_51_T_3[6:0] ? myVec_80 : _GEN_9977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9979 = 7'h51 == _myNewVec_51_T_3[6:0] ? myVec_81 : _GEN_9978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9980 = 7'h52 == _myNewVec_51_T_3[6:0] ? myVec_82 : _GEN_9979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9981 = 7'h53 == _myNewVec_51_T_3[6:0] ? myVec_83 : _GEN_9980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9982 = 7'h54 == _myNewVec_51_T_3[6:0] ? myVec_84 : _GEN_9981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9983 = 7'h55 == _myNewVec_51_T_3[6:0] ? myVec_85 : _GEN_9982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9984 = 7'h56 == _myNewVec_51_T_3[6:0] ? myVec_86 : _GEN_9983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9985 = 7'h57 == _myNewVec_51_T_3[6:0] ? myVec_87 : _GEN_9984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9986 = 7'h58 == _myNewVec_51_T_3[6:0] ? myVec_88 : _GEN_9985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9987 = 7'h59 == _myNewVec_51_T_3[6:0] ? myVec_89 : _GEN_9986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9988 = 7'h5a == _myNewVec_51_T_3[6:0] ? myVec_90 : _GEN_9987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9989 = 7'h5b == _myNewVec_51_T_3[6:0] ? myVec_91 : _GEN_9988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9990 = 7'h5c == _myNewVec_51_T_3[6:0] ? myVec_92 : _GEN_9989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9991 = 7'h5d == _myNewVec_51_T_3[6:0] ? myVec_93 : _GEN_9990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9992 = 7'h5e == _myNewVec_51_T_3[6:0] ? myVec_94 : _GEN_9991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9993 = 7'h5f == _myNewVec_51_T_3[6:0] ? myVec_95 : _GEN_9992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9994 = 7'h60 == _myNewVec_51_T_3[6:0] ? myVec_96 : _GEN_9993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9995 = 7'h61 == _myNewVec_51_T_3[6:0] ? myVec_97 : _GEN_9994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9996 = 7'h62 == _myNewVec_51_T_3[6:0] ? myVec_98 : _GEN_9995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9997 = 7'h63 == _myNewVec_51_T_3[6:0] ? myVec_99 : _GEN_9996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9998 = 7'h64 == _myNewVec_51_T_3[6:0] ? myVec_100 : _GEN_9997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_9999 = 7'h65 == _myNewVec_51_T_3[6:0] ? myVec_101 : _GEN_9998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10000 = 7'h66 == _myNewVec_51_T_3[6:0] ? myVec_102 : _GEN_9999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10001 = 7'h67 == _myNewVec_51_T_3[6:0] ? myVec_103 : _GEN_10000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10002 = 7'h68 == _myNewVec_51_T_3[6:0] ? myVec_104 : _GEN_10001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10003 = 7'h69 == _myNewVec_51_T_3[6:0] ? myVec_105 : _GEN_10002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10004 = 7'h6a == _myNewVec_51_T_3[6:0] ? myVec_106 : _GEN_10003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10005 = 7'h6b == _myNewVec_51_T_3[6:0] ? myVec_107 : _GEN_10004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10006 = 7'h6c == _myNewVec_51_T_3[6:0] ? myVec_108 : _GEN_10005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10007 = 7'h6d == _myNewVec_51_T_3[6:0] ? myVec_109 : _GEN_10006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10008 = 7'h6e == _myNewVec_51_T_3[6:0] ? myVec_110 : _GEN_10007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10009 = 7'h6f == _myNewVec_51_T_3[6:0] ? myVec_111 : _GEN_10008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10010 = 7'h70 == _myNewVec_51_T_3[6:0] ? myVec_112 : _GEN_10009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10011 = 7'h71 == _myNewVec_51_T_3[6:0] ? myVec_113 : _GEN_10010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10012 = 7'h72 == _myNewVec_51_T_3[6:0] ? myVec_114 : _GEN_10011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10013 = 7'h73 == _myNewVec_51_T_3[6:0] ? myVec_115 : _GEN_10012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10014 = 7'h74 == _myNewVec_51_T_3[6:0] ? myVec_116 : _GEN_10013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10015 = 7'h75 == _myNewVec_51_T_3[6:0] ? myVec_117 : _GEN_10014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10016 = 7'h76 == _myNewVec_51_T_3[6:0] ? myVec_118 : _GEN_10015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10017 = 7'h77 == _myNewVec_51_T_3[6:0] ? myVec_119 : _GEN_10016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10018 = 7'h78 == _myNewVec_51_T_3[6:0] ? myVec_120 : _GEN_10017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10019 = 7'h79 == _myNewVec_51_T_3[6:0] ? myVec_121 : _GEN_10018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10020 = 7'h7a == _myNewVec_51_T_3[6:0] ? myVec_122 : _GEN_10019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10021 = 7'h7b == _myNewVec_51_T_3[6:0] ? myVec_123 : _GEN_10020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10022 = 7'h7c == _myNewVec_51_T_3[6:0] ? myVec_124 : _GEN_10021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10023 = 7'h7d == _myNewVec_51_T_3[6:0] ? myVec_125 : _GEN_10022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10024 = 7'h7e == _myNewVec_51_T_3[6:0] ? myVec_126 : _GEN_10023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_51 = 7'h7f == _myNewVec_51_T_3[6:0] ? myVec_127 : _GEN_10024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_50_T_3 = _myNewVec_127_T_1 + 16'h4d; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_10027 = 7'h1 == _myNewVec_50_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10028 = 7'h2 == _myNewVec_50_T_3[6:0] ? myVec_2 : _GEN_10027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10029 = 7'h3 == _myNewVec_50_T_3[6:0] ? myVec_3 : _GEN_10028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10030 = 7'h4 == _myNewVec_50_T_3[6:0] ? myVec_4 : _GEN_10029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10031 = 7'h5 == _myNewVec_50_T_3[6:0] ? myVec_5 : _GEN_10030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10032 = 7'h6 == _myNewVec_50_T_3[6:0] ? myVec_6 : _GEN_10031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10033 = 7'h7 == _myNewVec_50_T_3[6:0] ? myVec_7 : _GEN_10032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10034 = 7'h8 == _myNewVec_50_T_3[6:0] ? myVec_8 : _GEN_10033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10035 = 7'h9 == _myNewVec_50_T_3[6:0] ? myVec_9 : _GEN_10034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10036 = 7'ha == _myNewVec_50_T_3[6:0] ? myVec_10 : _GEN_10035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10037 = 7'hb == _myNewVec_50_T_3[6:0] ? myVec_11 : _GEN_10036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10038 = 7'hc == _myNewVec_50_T_3[6:0] ? myVec_12 : _GEN_10037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10039 = 7'hd == _myNewVec_50_T_3[6:0] ? myVec_13 : _GEN_10038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10040 = 7'he == _myNewVec_50_T_3[6:0] ? myVec_14 : _GEN_10039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10041 = 7'hf == _myNewVec_50_T_3[6:0] ? myVec_15 : _GEN_10040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10042 = 7'h10 == _myNewVec_50_T_3[6:0] ? myVec_16 : _GEN_10041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10043 = 7'h11 == _myNewVec_50_T_3[6:0] ? myVec_17 : _GEN_10042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10044 = 7'h12 == _myNewVec_50_T_3[6:0] ? myVec_18 : _GEN_10043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10045 = 7'h13 == _myNewVec_50_T_3[6:0] ? myVec_19 : _GEN_10044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10046 = 7'h14 == _myNewVec_50_T_3[6:0] ? myVec_20 : _GEN_10045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10047 = 7'h15 == _myNewVec_50_T_3[6:0] ? myVec_21 : _GEN_10046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10048 = 7'h16 == _myNewVec_50_T_3[6:0] ? myVec_22 : _GEN_10047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10049 = 7'h17 == _myNewVec_50_T_3[6:0] ? myVec_23 : _GEN_10048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10050 = 7'h18 == _myNewVec_50_T_3[6:0] ? myVec_24 : _GEN_10049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10051 = 7'h19 == _myNewVec_50_T_3[6:0] ? myVec_25 : _GEN_10050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10052 = 7'h1a == _myNewVec_50_T_3[6:0] ? myVec_26 : _GEN_10051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10053 = 7'h1b == _myNewVec_50_T_3[6:0] ? myVec_27 : _GEN_10052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10054 = 7'h1c == _myNewVec_50_T_3[6:0] ? myVec_28 : _GEN_10053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10055 = 7'h1d == _myNewVec_50_T_3[6:0] ? myVec_29 : _GEN_10054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10056 = 7'h1e == _myNewVec_50_T_3[6:0] ? myVec_30 : _GEN_10055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10057 = 7'h1f == _myNewVec_50_T_3[6:0] ? myVec_31 : _GEN_10056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10058 = 7'h20 == _myNewVec_50_T_3[6:0] ? myVec_32 : _GEN_10057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10059 = 7'h21 == _myNewVec_50_T_3[6:0] ? myVec_33 : _GEN_10058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10060 = 7'h22 == _myNewVec_50_T_3[6:0] ? myVec_34 : _GEN_10059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10061 = 7'h23 == _myNewVec_50_T_3[6:0] ? myVec_35 : _GEN_10060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10062 = 7'h24 == _myNewVec_50_T_3[6:0] ? myVec_36 : _GEN_10061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10063 = 7'h25 == _myNewVec_50_T_3[6:0] ? myVec_37 : _GEN_10062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10064 = 7'h26 == _myNewVec_50_T_3[6:0] ? myVec_38 : _GEN_10063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10065 = 7'h27 == _myNewVec_50_T_3[6:0] ? myVec_39 : _GEN_10064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10066 = 7'h28 == _myNewVec_50_T_3[6:0] ? myVec_40 : _GEN_10065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10067 = 7'h29 == _myNewVec_50_T_3[6:0] ? myVec_41 : _GEN_10066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10068 = 7'h2a == _myNewVec_50_T_3[6:0] ? myVec_42 : _GEN_10067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10069 = 7'h2b == _myNewVec_50_T_3[6:0] ? myVec_43 : _GEN_10068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10070 = 7'h2c == _myNewVec_50_T_3[6:0] ? myVec_44 : _GEN_10069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10071 = 7'h2d == _myNewVec_50_T_3[6:0] ? myVec_45 : _GEN_10070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10072 = 7'h2e == _myNewVec_50_T_3[6:0] ? myVec_46 : _GEN_10071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10073 = 7'h2f == _myNewVec_50_T_3[6:0] ? myVec_47 : _GEN_10072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10074 = 7'h30 == _myNewVec_50_T_3[6:0] ? myVec_48 : _GEN_10073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10075 = 7'h31 == _myNewVec_50_T_3[6:0] ? myVec_49 : _GEN_10074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10076 = 7'h32 == _myNewVec_50_T_3[6:0] ? myVec_50 : _GEN_10075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10077 = 7'h33 == _myNewVec_50_T_3[6:0] ? myVec_51 : _GEN_10076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10078 = 7'h34 == _myNewVec_50_T_3[6:0] ? myVec_52 : _GEN_10077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10079 = 7'h35 == _myNewVec_50_T_3[6:0] ? myVec_53 : _GEN_10078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10080 = 7'h36 == _myNewVec_50_T_3[6:0] ? myVec_54 : _GEN_10079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10081 = 7'h37 == _myNewVec_50_T_3[6:0] ? myVec_55 : _GEN_10080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10082 = 7'h38 == _myNewVec_50_T_3[6:0] ? myVec_56 : _GEN_10081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10083 = 7'h39 == _myNewVec_50_T_3[6:0] ? myVec_57 : _GEN_10082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10084 = 7'h3a == _myNewVec_50_T_3[6:0] ? myVec_58 : _GEN_10083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10085 = 7'h3b == _myNewVec_50_T_3[6:0] ? myVec_59 : _GEN_10084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10086 = 7'h3c == _myNewVec_50_T_3[6:0] ? myVec_60 : _GEN_10085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10087 = 7'h3d == _myNewVec_50_T_3[6:0] ? myVec_61 : _GEN_10086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10088 = 7'h3e == _myNewVec_50_T_3[6:0] ? myVec_62 : _GEN_10087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10089 = 7'h3f == _myNewVec_50_T_3[6:0] ? myVec_63 : _GEN_10088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10090 = 7'h40 == _myNewVec_50_T_3[6:0] ? myVec_64 : _GEN_10089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10091 = 7'h41 == _myNewVec_50_T_3[6:0] ? myVec_65 : _GEN_10090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10092 = 7'h42 == _myNewVec_50_T_3[6:0] ? myVec_66 : _GEN_10091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10093 = 7'h43 == _myNewVec_50_T_3[6:0] ? myVec_67 : _GEN_10092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10094 = 7'h44 == _myNewVec_50_T_3[6:0] ? myVec_68 : _GEN_10093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10095 = 7'h45 == _myNewVec_50_T_3[6:0] ? myVec_69 : _GEN_10094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10096 = 7'h46 == _myNewVec_50_T_3[6:0] ? myVec_70 : _GEN_10095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10097 = 7'h47 == _myNewVec_50_T_3[6:0] ? myVec_71 : _GEN_10096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10098 = 7'h48 == _myNewVec_50_T_3[6:0] ? myVec_72 : _GEN_10097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10099 = 7'h49 == _myNewVec_50_T_3[6:0] ? myVec_73 : _GEN_10098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10100 = 7'h4a == _myNewVec_50_T_3[6:0] ? myVec_74 : _GEN_10099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10101 = 7'h4b == _myNewVec_50_T_3[6:0] ? myVec_75 : _GEN_10100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10102 = 7'h4c == _myNewVec_50_T_3[6:0] ? myVec_76 : _GEN_10101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10103 = 7'h4d == _myNewVec_50_T_3[6:0] ? myVec_77 : _GEN_10102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10104 = 7'h4e == _myNewVec_50_T_3[6:0] ? myVec_78 : _GEN_10103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10105 = 7'h4f == _myNewVec_50_T_3[6:0] ? myVec_79 : _GEN_10104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10106 = 7'h50 == _myNewVec_50_T_3[6:0] ? myVec_80 : _GEN_10105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10107 = 7'h51 == _myNewVec_50_T_3[6:0] ? myVec_81 : _GEN_10106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10108 = 7'h52 == _myNewVec_50_T_3[6:0] ? myVec_82 : _GEN_10107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10109 = 7'h53 == _myNewVec_50_T_3[6:0] ? myVec_83 : _GEN_10108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10110 = 7'h54 == _myNewVec_50_T_3[6:0] ? myVec_84 : _GEN_10109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10111 = 7'h55 == _myNewVec_50_T_3[6:0] ? myVec_85 : _GEN_10110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10112 = 7'h56 == _myNewVec_50_T_3[6:0] ? myVec_86 : _GEN_10111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10113 = 7'h57 == _myNewVec_50_T_3[6:0] ? myVec_87 : _GEN_10112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10114 = 7'h58 == _myNewVec_50_T_3[6:0] ? myVec_88 : _GEN_10113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10115 = 7'h59 == _myNewVec_50_T_3[6:0] ? myVec_89 : _GEN_10114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10116 = 7'h5a == _myNewVec_50_T_3[6:0] ? myVec_90 : _GEN_10115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10117 = 7'h5b == _myNewVec_50_T_3[6:0] ? myVec_91 : _GEN_10116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10118 = 7'h5c == _myNewVec_50_T_3[6:0] ? myVec_92 : _GEN_10117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10119 = 7'h5d == _myNewVec_50_T_3[6:0] ? myVec_93 : _GEN_10118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10120 = 7'h5e == _myNewVec_50_T_3[6:0] ? myVec_94 : _GEN_10119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10121 = 7'h5f == _myNewVec_50_T_3[6:0] ? myVec_95 : _GEN_10120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10122 = 7'h60 == _myNewVec_50_T_3[6:0] ? myVec_96 : _GEN_10121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10123 = 7'h61 == _myNewVec_50_T_3[6:0] ? myVec_97 : _GEN_10122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10124 = 7'h62 == _myNewVec_50_T_3[6:0] ? myVec_98 : _GEN_10123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10125 = 7'h63 == _myNewVec_50_T_3[6:0] ? myVec_99 : _GEN_10124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10126 = 7'h64 == _myNewVec_50_T_3[6:0] ? myVec_100 : _GEN_10125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10127 = 7'h65 == _myNewVec_50_T_3[6:0] ? myVec_101 : _GEN_10126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10128 = 7'h66 == _myNewVec_50_T_3[6:0] ? myVec_102 : _GEN_10127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10129 = 7'h67 == _myNewVec_50_T_3[6:0] ? myVec_103 : _GEN_10128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10130 = 7'h68 == _myNewVec_50_T_3[6:0] ? myVec_104 : _GEN_10129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10131 = 7'h69 == _myNewVec_50_T_3[6:0] ? myVec_105 : _GEN_10130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10132 = 7'h6a == _myNewVec_50_T_3[6:0] ? myVec_106 : _GEN_10131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10133 = 7'h6b == _myNewVec_50_T_3[6:0] ? myVec_107 : _GEN_10132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10134 = 7'h6c == _myNewVec_50_T_3[6:0] ? myVec_108 : _GEN_10133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10135 = 7'h6d == _myNewVec_50_T_3[6:0] ? myVec_109 : _GEN_10134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10136 = 7'h6e == _myNewVec_50_T_3[6:0] ? myVec_110 : _GEN_10135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10137 = 7'h6f == _myNewVec_50_T_3[6:0] ? myVec_111 : _GEN_10136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10138 = 7'h70 == _myNewVec_50_T_3[6:0] ? myVec_112 : _GEN_10137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10139 = 7'h71 == _myNewVec_50_T_3[6:0] ? myVec_113 : _GEN_10138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10140 = 7'h72 == _myNewVec_50_T_3[6:0] ? myVec_114 : _GEN_10139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10141 = 7'h73 == _myNewVec_50_T_3[6:0] ? myVec_115 : _GEN_10140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10142 = 7'h74 == _myNewVec_50_T_3[6:0] ? myVec_116 : _GEN_10141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10143 = 7'h75 == _myNewVec_50_T_3[6:0] ? myVec_117 : _GEN_10142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10144 = 7'h76 == _myNewVec_50_T_3[6:0] ? myVec_118 : _GEN_10143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10145 = 7'h77 == _myNewVec_50_T_3[6:0] ? myVec_119 : _GEN_10144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10146 = 7'h78 == _myNewVec_50_T_3[6:0] ? myVec_120 : _GEN_10145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10147 = 7'h79 == _myNewVec_50_T_3[6:0] ? myVec_121 : _GEN_10146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10148 = 7'h7a == _myNewVec_50_T_3[6:0] ? myVec_122 : _GEN_10147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10149 = 7'h7b == _myNewVec_50_T_3[6:0] ? myVec_123 : _GEN_10148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10150 = 7'h7c == _myNewVec_50_T_3[6:0] ? myVec_124 : _GEN_10149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10151 = 7'h7d == _myNewVec_50_T_3[6:0] ? myVec_125 : _GEN_10150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10152 = 7'h7e == _myNewVec_50_T_3[6:0] ? myVec_126 : _GEN_10151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_50 = 7'h7f == _myNewVec_50_T_3[6:0] ? myVec_127 : _GEN_10152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_49_T_3 = _myNewVec_127_T_1 + 16'h4e; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_10155 = 7'h1 == _myNewVec_49_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10156 = 7'h2 == _myNewVec_49_T_3[6:0] ? myVec_2 : _GEN_10155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10157 = 7'h3 == _myNewVec_49_T_3[6:0] ? myVec_3 : _GEN_10156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10158 = 7'h4 == _myNewVec_49_T_3[6:0] ? myVec_4 : _GEN_10157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10159 = 7'h5 == _myNewVec_49_T_3[6:0] ? myVec_5 : _GEN_10158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10160 = 7'h6 == _myNewVec_49_T_3[6:0] ? myVec_6 : _GEN_10159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10161 = 7'h7 == _myNewVec_49_T_3[6:0] ? myVec_7 : _GEN_10160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10162 = 7'h8 == _myNewVec_49_T_3[6:0] ? myVec_8 : _GEN_10161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10163 = 7'h9 == _myNewVec_49_T_3[6:0] ? myVec_9 : _GEN_10162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10164 = 7'ha == _myNewVec_49_T_3[6:0] ? myVec_10 : _GEN_10163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10165 = 7'hb == _myNewVec_49_T_3[6:0] ? myVec_11 : _GEN_10164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10166 = 7'hc == _myNewVec_49_T_3[6:0] ? myVec_12 : _GEN_10165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10167 = 7'hd == _myNewVec_49_T_3[6:0] ? myVec_13 : _GEN_10166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10168 = 7'he == _myNewVec_49_T_3[6:0] ? myVec_14 : _GEN_10167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10169 = 7'hf == _myNewVec_49_T_3[6:0] ? myVec_15 : _GEN_10168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10170 = 7'h10 == _myNewVec_49_T_3[6:0] ? myVec_16 : _GEN_10169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10171 = 7'h11 == _myNewVec_49_T_3[6:0] ? myVec_17 : _GEN_10170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10172 = 7'h12 == _myNewVec_49_T_3[6:0] ? myVec_18 : _GEN_10171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10173 = 7'h13 == _myNewVec_49_T_3[6:0] ? myVec_19 : _GEN_10172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10174 = 7'h14 == _myNewVec_49_T_3[6:0] ? myVec_20 : _GEN_10173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10175 = 7'h15 == _myNewVec_49_T_3[6:0] ? myVec_21 : _GEN_10174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10176 = 7'h16 == _myNewVec_49_T_3[6:0] ? myVec_22 : _GEN_10175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10177 = 7'h17 == _myNewVec_49_T_3[6:0] ? myVec_23 : _GEN_10176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10178 = 7'h18 == _myNewVec_49_T_3[6:0] ? myVec_24 : _GEN_10177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10179 = 7'h19 == _myNewVec_49_T_3[6:0] ? myVec_25 : _GEN_10178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10180 = 7'h1a == _myNewVec_49_T_3[6:0] ? myVec_26 : _GEN_10179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10181 = 7'h1b == _myNewVec_49_T_3[6:0] ? myVec_27 : _GEN_10180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10182 = 7'h1c == _myNewVec_49_T_3[6:0] ? myVec_28 : _GEN_10181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10183 = 7'h1d == _myNewVec_49_T_3[6:0] ? myVec_29 : _GEN_10182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10184 = 7'h1e == _myNewVec_49_T_3[6:0] ? myVec_30 : _GEN_10183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10185 = 7'h1f == _myNewVec_49_T_3[6:0] ? myVec_31 : _GEN_10184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10186 = 7'h20 == _myNewVec_49_T_3[6:0] ? myVec_32 : _GEN_10185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10187 = 7'h21 == _myNewVec_49_T_3[6:0] ? myVec_33 : _GEN_10186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10188 = 7'h22 == _myNewVec_49_T_3[6:0] ? myVec_34 : _GEN_10187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10189 = 7'h23 == _myNewVec_49_T_3[6:0] ? myVec_35 : _GEN_10188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10190 = 7'h24 == _myNewVec_49_T_3[6:0] ? myVec_36 : _GEN_10189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10191 = 7'h25 == _myNewVec_49_T_3[6:0] ? myVec_37 : _GEN_10190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10192 = 7'h26 == _myNewVec_49_T_3[6:0] ? myVec_38 : _GEN_10191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10193 = 7'h27 == _myNewVec_49_T_3[6:0] ? myVec_39 : _GEN_10192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10194 = 7'h28 == _myNewVec_49_T_3[6:0] ? myVec_40 : _GEN_10193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10195 = 7'h29 == _myNewVec_49_T_3[6:0] ? myVec_41 : _GEN_10194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10196 = 7'h2a == _myNewVec_49_T_3[6:0] ? myVec_42 : _GEN_10195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10197 = 7'h2b == _myNewVec_49_T_3[6:0] ? myVec_43 : _GEN_10196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10198 = 7'h2c == _myNewVec_49_T_3[6:0] ? myVec_44 : _GEN_10197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10199 = 7'h2d == _myNewVec_49_T_3[6:0] ? myVec_45 : _GEN_10198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10200 = 7'h2e == _myNewVec_49_T_3[6:0] ? myVec_46 : _GEN_10199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10201 = 7'h2f == _myNewVec_49_T_3[6:0] ? myVec_47 : _GEN_10200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10202 = 7'h30 == _myNewVec_49_T_3[6:0] ? myVec_48 : _GEN_10201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10203 = 7'h31 == _myNewVec_49_T_3[6:0] ? myVec_49 : _GEN_10202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10204 = 7'h32 == _myNewVec_49_T_3[6:0] ? myVec_50 : _GEN_10203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10205 = 7'h33 == _myNewVec_49_T_3[6:0] ? myVec_51 : _GEN_10204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10206 = 7'h34 == _myNewVec_49_T_3[6:0] ? myVec_52 : _GEN_10205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10207 = 7'h35 == _myNewVec_49_T_3[6:0] ? myVec_53 : _GEN_10206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10208 = 7'h36 == _myNewVec_49_T_3[6:0] ? myVec_54 : _GEN_10207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10209 = 7'h37 == _myNewVec_49_T_3[6:0] ? myVec_55 : _GEN_10208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10210 = 7'h38 == _myNewVec_49_T_3[6:0] ? myVec_56 : _GEN_10209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10211 = 7'h39 == _myNewVec_49_T_3[6:0] ? myVec_57 : _GEN_10210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10212 = 7'h3a == _myNewVec_49_T_3[6:0] ? myVec_58 : _GEN_10211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10213 = 7'h3b == _myNewVec_49_T_3[6:0] ? myVec_59 : _GEN_10212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10214 = 7'h3c == _myNewVec_49_T_3[6:0] ? myVec_60 : _GEN_10213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10215 = 7'h3d == _myNewVec_49_T_3[6:0] ? myVec_61 : _GEN_10214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10216 = 7'h3e == _myNewVec_49_T_3[6:0] ? myVec_62 : _GEN_10215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10217 = 7'h3f == _myNewVec_49_T_3[6:0] ? myVec_63 : _GEN_10216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10218 = 7'h40 == _myNewVec_49_T_3[6:0] ? myVec_64 : _GEN_10217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10219 = 7'h41 == _myNewVec_49_T_3[6:0] ? myVec_65 : _GEN_10218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10220 = 7'h42 == _myNewVec_49_T_3[6:0] ? myVec_66 : _GEN_10219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10221 = 7'h43 == _myNewVec_49_T_3[6:0] ? myVec_67 : _GEN_10220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10222 = 7'h44 == _myNewVec_49_T_3[6:0] ? myVec_68 : _GEN_10221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10223 = 7'h45 == _myNewVec_49_T_3[6:0] ? myVec_69 : _GEN_10222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10224 = 7'h46 == _myNewVec_49_T_3[6:0] ? myVec_70 : _GEN_10223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10225 = 7'h47 == _myNewVec_49_T_3[6:0] ? myVec_71 : _GEN_10224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10226 = 7'h48 == _myNewVec_49_T_3[6:0] ? myVec_72 : _GEN_10225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10227 = 7'h49 == _myNewVec_49_T_3[6:0] ? myVec_73 : _GEN_10226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10228 = 7'h4a == _myNewVec_49_T_3[6:0] ? myVec_74 : _GEN_10227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10229 = 7'h4b == _myNewVec_49_T_3[6:0] ? myVec_75 : _GEN_10228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10230 = 7'h4c == _myNewVec_49_T_3[6:0] ? myVec_76 : _GEN_10229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10231 = 7'h4d == _myNewVec_49_T_3[6:0] ? myVec_77 : _GEN_10230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10232 = 7'h4e == _myNewVec_49_T_3[6:0] ? myVec_78 : _GEN_10231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10233 = 7'h4f == _myNewVec_49_T_3[6:0] ? myVec_79 : _GEN_10232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10234 = 7'h50 == _myNewVec_49_T_3[6:0] ? myVec_80 : _GEN_10233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10235 = 7'h51 == _myNewVec_49_T_3[6:0] ? myVec_81 : _GEN_10234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10236 = 7'h52 == _myNewVec_49_T_3[6:0] ? myVec_82 : _GEN_10235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10237 = 7'h53 == _myNewVec_49_T_3[6:0] ? myVec_83 : _GEN_10236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10238 = 7'h54 == _myNewVec_49_T_3[6:0] ? myVec_84 : _GEN_10237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10239 = 7'h55 == _myNewVec_49_T_3[6:0] ? myVec_85 : _GEN_10238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10240 = 7'h56 == _myNewVec_49_T_3[6:0] ? myVec_86 : _GEN_10239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10241 = 7'h57 == _myNewVec_49_T_3[6:0] ? myVec_87 : _GEN_10240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10242 = 7'h58 == _myNewVec_49_T_3[6:0] ? myVec_88 : _GEN_10241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10243 = 7'h59 == _myNewVec_49_T_3[6:0] ? myVec_89 : _GEN_10242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10244 = 7'h5a == _myNewVec_49_T_3[6:0] ? myVec_90 : _GEN_10243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10245 = 7'h5b == _myNewVec_49_T_3[6:0] ? myVec_91 : _GEN_10244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10246 = 7'h5c == _myNewVec_49_T_3[6:0] ? myVec_92 : _GEN_10245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10247 = 7'h5d == _myNewVec_49_T_3[6:0] ? myVec_93 : _GEN_10246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10248 = 7'h5e == _myNewVec_49_T_3[6:0] ? myVec_94 : _GEN_10247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10249 = 7'h5f == _myNewVec_49_T_3[6:0] ? myVec_95 : _GEN_10248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10250 = 7'h60 == _myNewVec_49_T_3[6:0] ? myVec_96 : _GEN_10249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10251 = 7'h61 == _myNewVec_49_T_3[6:0] ? myVec_97 : _GEN_10250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10252 = 7'h62 == _myNewVec_49_T_3[6:0] ? myVec_98 : _GEN_10251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10253 = 7'h63 == _myNewVec_49_T_3[6:0] ? myVec_99 : _GEN_10252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10254 = 7'h64 == _myNewVec_49_T_3[6:0] ? myVec_100 : _GEN_10253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10255 = 7'h65 == _myNewVec_49_T_3[6:0] ? myVec_101 : _GEN_10254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10256 = 7'h66 == _myNewVec_49_T_3[6:0] ? myVec_102 : _GEN_10255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10257 = 7'h67 == _myNewVec_49_T_3[6:0] ? myVec_103 : _GEN_10256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10258 = 7'h68 == _myNewVec_49_T_3[6:0] ? myVec_104 : _GEN_10257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10259 = 7'h69 == _myNewVec_49_T_3[6:0] ? myVec_105 : _GEN_10258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10260 = 7'h6a == _myNewVec_49_T_3[6:0] ? myVec_106 : _GEN_10259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10261 = 7'h6b == _myNewVec_49_T_3[6:0] ? myVec_107 : _GEN_10260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10262 = 7'h6c == _myNewVec_49_T_3[6:0] ? myVec_108 : _GEN_10261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10263 = 7'h6d == _myNewVec_49_T_3[6:0] ? myVec_109 : _GEN_10262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10264 = 7'h6e == _myNewVec_49_T_3[6:0] ? myVec_110 : _GEN_10263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10265 = 7'h6f == _myNewVec_49_T_3[6:0] ? myVec_111 : _GEN_10264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10266 = 7'h70 == _myNewVec_49_T_3[6:0] ? myVec_112 : _GEN_10265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10267 = 7'h71 == _myNewVec_49_T_3[6:0] ? myVec_113 : _GEN_10266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10268 = 7'h72 == _myNewVec_49_T_3[6:0] ? myVec_114 : _GEN_10267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10269 = 7'h73 == _myNewVec_49_T_3[6:0] ? myVec_115 : _GEN_10268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10270 = 7'h74 == _myNewVec_49_T_3[6:0] ? myVec_116 : _GEN_10269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10271 = 7'h75 == _myNewVec_49_T_3[6:0] ? myVec_117 : _GEN_10270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10272 = 7'h76 == _myNewVec_49_T_3[6:0] ? myVec_118 : _GEN_10271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10273 = 7'h77 == _myNewVec_49_T_3[6:0] ? myVec_119 : _GEN_10272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10274 = 7'h78 == _myNewVec_49_T_3[6:0] ? myVec_120 : _GEN_10273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10275 = 7'h79 == _myNewVec_49_T_3[6:0] ? myVec_121 : _GEN_10274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10276 = 7'h7a == _myNewVec_49_T_3[6:0] ? myVec_122 : _GEN_10275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10277 = 7'h7b == _myNewVec_49_T_3[6:0] ? myVec_123 : _GEN_10276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10278 = 7'h7c == _myNewVec_49_T_3[6:0] ? myVec_124 : _GEN_10277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10279 = 7'h7d == _myNewVec_49_T_3[6:0] ? myVec_125 : _GEN_10278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10280 = 7'h7e == _myNewVec_49_T_3[6:0] ? myVec_126 : _GEN_10279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_49 = 7'h7f == _myNewVec_49_T_3[6:0] ? myVec_127 : _GEN_10280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_48_T_3 = _myNewVec_127_T_1 + 16'h4f; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_10283 = 7'h1 == _myNewVec_48_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10284 = 7'h2 == _myNewVec_48_T_3[6:0] ? myVec_2 : _GEN_10283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10285 = 7'h3 == _myNewVec_48_T_3[6:0] ? myVec_3 : _GEN_10284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10286 = 7'h4 == _myNewVec_48_T_3[6:0] ? myVec_4 : _GEN_10285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10287 = 7'h5 == _myNewVec_48_T_3[6:0] ? myVec_5 : _GEN_10286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10288 = 7'h6 == _myNewVec_48_T_3[6:0] ? myVec_6 : _GEN_10287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10289 = 7'h7 == _myNewVec_48_T_3[6:0] ? myVec_7 : _GEN_10288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10290 = 7'h8 == _myNewVec_48_T_3[6:0] ? myVec_8 : _GEN_10289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10291 = 7'h9 == _myNewVec_48_T_3[6:0] ? myVec_9 : _GEN_10290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10292 = 7'ha == _myNewVec_48_T_3[6:0] ? myVec_10 : _GEN_10291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10293 = 7'hb == _myNewVec_48_T_3[6:0] ? myVec_11 : _GEN_10292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10294 = 7'hc == _myNewVec_48_T_3[6:0] ? myVec_12 : _GEN_10293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10295 = 7'hd == _myNewVec_48_T_3[6:0] ? myVec_13 : _GEN_10294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10296 = 7'he == _myNewVec_48_T_3[6:0] ? myVec_14 : _GEN_10295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10297 = 7'hf == _myNewVec_48_T_3[6:0] ? myVec_15 : _GEN_10296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10298 = 7'h10 == _myNewVec_48_T_3[6:0] ? myVec_16 : _GEN_10297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10299 = 7'h11 == _myNewVec_48_T_3[6:0] ? myVec_17 : _GEN_10298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10300 = 7'h12 == _myNewVec_48_T_3[6:0] ? myVec_18 : _GEN_10299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10301 = 7'h13 == _myNewVec_48_T_3[6:0] ? myVec_19 : _GEN_10300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10302 = 7'h14 == _myNewVec_48_T_3[6:0] ? myVec_20 : _GEN_10301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10303 = 7'h15 == _myNewVec_48_T_3[6:0] ? myVec_21 : _GEN_10302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10304 = 7'h16 == _myNewVec_48_T_3[6:0] ? myVec_22 : _GEN_10303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10305 = 7'h17 == _myNewVec_48_T_3[6:0] ? myVec_23 : _GEN_10304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10306 = 7'h18 == _myNewVec_48_T_3[6:0] ? myVec_24 : _GEN_10305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10307 = 7'h19 == _myNewVec_48_T_3[6:0] ? myVec_25 : _GEN_10306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10308 = 7'h1a == _myNewVec_48_T_3[6:0] ? myVec_26 : _GEN_10307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10309 = 7'h1b == _myNewVec_48_T_3[6:0] ? myVec_27 : _GEN_10308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10310 = 7'h1c == _myNewVec_48_T_3[6:0] ? myVec_28 : _GEN_10309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10311 = 7'h1d == _myNewVec_48_T_3[6:0] ? myVec_29 : _GEN_10310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10312 = 7'h1e == _myNewVec_48_T_3[6:0] ? myVec_30 : _GEN_10311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10313 = 7'h1f == _myNewVec_48_T_3[6:0] ? myVec_31 : _GEN_10312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10314 = 7'h20 == _myNewVec_48_T_3[6:0] ? myVec_32 : _GEN_10313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10315 = 7'h21 == _myNewVec_48_T_3[6:0] ? myVec_33 : _GEN_10314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10316 = 7'h22 == _myNewVec_48_T_3[6:0] ? myVec_34 : _GEN_10315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10317 = 7'h23 == _myNewVec_48_T_3[6:0] ? myVec_35 : _GEN_10316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10318 = 7'h24 == _myNewVec_48_T_3[6:0] ? myVec_36 : _GEN_10317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10319 = 7'h25 == _myNewVec_48_T_3[6:0] ? myVec_37 : _GEN_10318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10320 = 7'h26 == _myNewVec_48_T_3[6:0] ? myVec_38 : _GEN_10319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10321 = 7'h27 == _myNewVec_48_T_3[6:0] ? myVec_39 : _GEN_10320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10322 = 7'h28 == _myNewVec_48_T_3[6:0] ? myVec_40 : _GEN_10321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10323 = 7'h29 == _myNewVec_48_T_3[6:0] ? myVec_41 : _GEN_10322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10324 = 7'h2a == _myNewVec_48_T_3[6:0] ? myVec_42 : _GEN_10323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10325 = 7'h2b == _myNewVec_48_T_3[6:0] ? myVec_43 : _GEN_10324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10326 = 7'h2c == _myNewVec_48_T_3[6:0] ? myVec_44 : _GEN_10325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10327 = 7'h2d == _myNewVec_48_T_3[6:0] ? myVec_45 : _GEN_10326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10328 = 7'h2e == _myNewVec_48_T_3[6:0] ? myVec_46 : _GEN_10327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10329 = 7'h2f == _myNewVec_48_T_3[6:0] ? myVec_47 : _GEN_10328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10330 = 7'h30 == _myNewVec_48_T_3[6:0] ? myVec_48 : _GEN_10329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10331 = 7'h31 == _myNewVec_48_T_3[6:0] ? myVec_49 : _GEN_10330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10332 = 7'h32 == _myNewVec_48_T_3[6:0] ? myVec_50 : _GEN_10331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10333 = 7'h33 == _myNewVec_48_T_3[6:0] ? myVec_51 : _GEN_10332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10334 = 7'h34 == _myNewVec_48_T_3[6:0] ? myVec_52 : _GEN_10333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10335 = 7'h35 == _myNewVec_48_T_3[6:0] ? myVec_53 : _GEN_10334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10336 = 7'h36 == _myNewVec_48_T_3[6:0] ? myVec_54 : _GEN_10335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10337 = 7'h37 == _myNewVec_48_T_3[6:0] ? myVec_55 : _GEN_10336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10338 = 7'h38 == _myNewVec_48_T_3[6:0] ? myVec_56 : _GEN_10337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10339 = 7'h39 == _myNewVec_48_T_3[6:0] ? myVec_57 : _GEN_10338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10340 = 7'h3a == _myNewVec_48_T_3[6:0] ? myVec_58 : _GEN_10339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10341 = 7'h3b == _myNewVec_48_T_3[6:0] ? myVec_59 : _GEN_10340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10342 = 7'h3c == _myNewVec_48_T_3[6:0] ? myVec_60 : _GEN_10341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10343 = 7'h3d == _myNewVec_48_T_3[6:0] ? myVec_61 : _GEN_10342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10344 = 7'h3e == _myNewVec_48_T_3[6:0] ? myVec_62 : _GEN_10343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10345 = 7'h3f == _myNewVec_48_T_3[6:0] ? myVec_63 : _GEN_10344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10346 = 7'h40 == _myNewVec_48_T_3[6:0] ? myVec_64 : _GEN_10345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10347 = 7'h41 == _myNewVec_48_T_3[6:0] ? myVec_65 : _GEN_10346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10348 = 7'h42 == _myNewVec_48_T_3[6:0] ? myVec_66 : _GEN_10347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10349 = 7'h43 == _myNewVec_48_T_3[6:0] ? myVec_67 : _GEN_10348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10350 = 7'h44 == _myNewVec_48_T_3[6:0] ? myVec_68 : _GEN_10349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10351 = 7'h45 == _myNewVec_48_T_3[6:0] ? myVec_69 : _GEN_10350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10352 = 7'h46 == _myNewVec_48_T_3[6:0] ? myVec_70 : _GEN_10351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10353 = 7'h47 == _myNewVec_48_T_3[6:0] ? myVec_71 : _GEN_10352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10354 = 7'h48 == _myNewVec_48_T_3[6:0] ? myVec_72 : _GEN_10353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10355 = 7'h49 == _myNewVec_48_T_3[6:0] ? myVec_73 : _GEN_10354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10356 = 7'h4a == _myNewVec_48_T_3[6:0] ? myVec_74 : _GEN_10355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10357 = 7'h4b == _myNewVec_48_T_3[6:0] ? myVec_75 : _GEN_10356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10358 = 7'h4c == _myNewVec_48_T_3[6:0] ? myVec_76 : _GEN_10357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10359 = 7'h4d == _myNewVec_48_T_3[6:0] ? myVec_77 : _GEN_10358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10360 = 7'h4e == _myNewVec_48_T_3[6:0] ? myVec_78 : _GEN_10359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10361 = 7'h4f == _myNewVec_48_T_3[6:0] ? myVec_79 : _GEN_10360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10362 = 7'h50 == _myNewVec_48_T_3[6:0] ? myVec_80 : _GEN_10361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10363 = 7'h51 == _myNewVec_48_T_3[6:0] ? myVec_81 : _GEN_10362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10364 = 7'h52 == _myNewVec_48_T_3[6:0] ? myVec_82 : _GEN_10363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10365 = 7'h53 == _myNewVec_48_T_3[6:0] ? myVec_83 : _GEN_10364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10366 = 7'h54 == _myNewVec_48_T_3[6:0] ? myVec_84 : _GEN_10365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10367 = 7'h55 == _myNewVec_48_T_3[6:0] ? myVec_85 : _GEN_10366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10368 = 7'h56 == _myNewVec_48_T_3[6:0] ? myVec_86 : _GEN_10367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10369 = 7'h57 == _myNewVec_48_T_3[6:0] ? myVec_87 : _GEN_10368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10370 = 7'h58 == _myNewVec_48_T_3[6:0] ? myVec_88 : _GEN_10369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10371 = 7'h59 == _myNewVec_48_T_3[6:0] ? myVec_89 : _GEN_10370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10372 = 7'h5a == _myNewVec_48_T_3[6:0] ? myVec_90 : _GEN_10371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10373 = 7'h5b == _myNewVec_48_T_3[6:0] ? myVec_91 : _GEN_10372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10374 = 7'h5c == _myNewVec_48_T_3[6:0] ? myVec_92 : _GEN_10373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10375 = 7'h5d == _myNewVec_48_T_3[6:0] ? myVec_93 : _GEN_10374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10376 = 7'h5e == _myNewVec_48_T_3[6:0] ? myVec_94 : _GEN_10375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10377 = 7'h5f == _myNewVec_48_T_3[6:0] ? myVec_95 : _GEN_10376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10378 = 7'h60 == _myNewVec_48_T_3[6:0] ? myVec_96 : _GEN_10377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10379 = 7'h61 == _myNewVec_48_T_3[6:0] ? myVec_97 : _GEN_10378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10380 = 7'h62 == _myNewVec_48_T_3[6:0] ? myVec_98 : _GEN_10379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10381 = 7'h63 == _myNewVec_48_T_3[6:0] ? myVec_99 : _GEN_10380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10382 = 7'h64 == _myNewVec_48_T_3[6:0] ? myVec_100 : _GEN_10381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10383 = 7'h65 == _myNewVec_48_T_3[6:0] ? myVec_101 : _GEN_10382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10384 = 7'h66 == _myNewVec_48_T_3[6:0] ? myVec_102 : _GEN_10383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10385 = 7'h67 == _myNewVec_48_T_3[6:0] ? myVec_103 : _GEN_10384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10386 = 7'h68 == _myNewVec_48_T_3[6:0] ? myVec_104 : _GEN_10385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10387 = 7'h69 == _myNewVec_48_T_3[6:0] ? myVec_105 : _GEN_10386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10388 = 7'h6a == _myNewVec_48_T_3[6:0] ? myVec_106 : _GEN_10387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10389 = 7'h6b == _myNewVec_48_T_3[6:0] ? myVec_107 : _GEN_10388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10390 = 7'h6c == _myNewVec_48_T_3[6:0] ? myVec_108 : _GEN_10389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10391 = 7'h6d == _myNewVec_48_T_3[6:0] ? myVec_109 : _GEN_10390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10392 = 7'h6e == _myNewVec_48_T_3[6:0] ? myVec_110 : _GEN_10391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10393 = 7'h6f == _myNewVec_48_T_3[6:0] ? myVec_111 : _GEN_10392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10394 = 7'h70 == _myNewVec_48_T_3[6:0] ? myVec_112 : _GEN_10393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10395 = 7'h71 == _myNewVec_48_T_3[6:0] ? myVec_113 : _GEN_10394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10396 = 7'h72 == _myNewVec_48_T_3[6:0] ? myVec_114 : _GEN_10395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10397 = 7'h73 == _myNewVec_48_T_3[6:0] ? myVec_115 : _GEN_10396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10398 = 7'h74 == _myNewVec_48_T_3[6:0] ? myVec_116 : _GEN_10397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10399 = 7'h75 == _myNewVec_48_T_3[6:0] ? myVec_117 : _GEN_10398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10400 = 7'h76 == _myNewVec_48_T_3[6:0] ? myVec_118 : _GEN_10399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10401 = 7'h77 == _myNewVec_48_T_3[6:0] ? myVec_119 : _GEN_10400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10402 = 7'h78 == _myNewVec_48_T_3[6:0] ? myVec_120 : _GEN_10401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10403 = 7'h79 == _myNewVec_48_T_3[6:0] ? myVec_121 : _GEN_10402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10404 = 7'h7a == _myNewVec_48_T_3[6:0] ? myVec_122 : _GEN_10403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10405 = 7'h7b == _myNewVec_48_T_3[6:0] ? myVec_123 : _GEN_10404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10406 = 7'h7c == _myNewVec_48_T_3[6:0] ? myVec_124 : _GEN_10405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10407 = 7'h7d == _myNewVec_48_T_3[6:0] ? myVec_125 : _GEN_10406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10408 = 7'h7e == _myNewVec_48_T_3[6:0] ? myVec_126 : _GEN_10407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_48 = 7'h7f == _myNewVec_48_T_3[6:0] ? myVec_127 : _GEN_10408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [255:0] myNewWire_lo_hi_hi_lo = {myNewVec_55,myNewVec_54,myNewVec_53,myNewVec_52,myNewVec_51,myNewVec_50,
    myNewVec_49,myNewVec_48}; // @[hh_datapath_chisel.scala 238:27]
  wire [15:0] _myNewVec_47_T_3 = _myNewVec_127_T_1 + 16'h50; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_10411 = 7'h1 == _myNewVec_47_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10412 = 7'h2 == _myNewVec_47_T_3[6:0] ? myVec_2 : _GEN_10411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10413 = 7'h3 == _myNewVec_47_T_3[6:0] ? myVec_3 : _GEN_10412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10414 = 7'h4 == _myNewVec_47_T_3[6:0] ? myVec_4 : _GEN_10413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10415 = 7'h5 == _myNewVec_47_T_3[6:0] ? myVec_5 : _GEN_10414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10416 = 7'h6 == _myNewVec_47_T_3[6:0] ? myVec_6 : _GEN_10415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10417 = 7'h7 == _myNewVec_47_T_3[6:0] ? myVec_7 : _GEN_10416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10418 = 7'h8 == _myNewVec_47_T_3[6:0] ? myVec_8 : _GEN_10417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10419 = 7'h9 == _myNewVec_47_T_3[6:0] ? myVec_9 : _GEN_10418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10420 = 7'ha == _myNewVec_47_T_3[6:0] ? myVec_10 : _GEN_10419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10421 = 7'hb == _myNewVec_47_T_3[6:0] ? myVec_11 : _GEN_10420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10422 = 7'hc == _myNewVec_47_T_3[6:0] ? myVec_12 : _GEN_10421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10423 = 7'hd == _myNewVec_47_T_3[6:0] ? myVec_13 : _GEN_10422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10424 = 7'he == _myNewVec_47_T_3[6:0] ? myVec_14 : _GEN_10423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10425 = 7'hf == _myNewVec_47_T_3[6:0] ? myVec_15 : _GEN_10424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10426 = 7'h10 == _myNewVec_47_T_3[6:0] ? myVec_16 : _GEN_10425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10427 = 7'h11 == _myNewVec_47_T_3[6:0] ? myVec_17 : _GEN_10426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10428 = 7'h12 == _myNewVec_47_T_3[6:0] ? myVec_18 : _GEN_10427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10429 = 7'h13 == _myNewVec_47_T_3[6:0] ? myVec_19 : _GEN_10428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10430 = 7'h14 == _myNewVec_47_T_3[6:0] ? myVec_20 : _GEN_10429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10431 = 7'h15 == _myNewVec_47_T_3[6:0] ? myVec_21 : _GEN_10430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10432 = 7'h16 == _myNewVec_47_T_3[6:0] ? myVec_22 : _GEN_10431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10433 = 7'h17 == _myNewVec_47_T_3[6:0] ? myVec_23 : _GEN_10432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10434 = 7'h18 == _myNewVec_47_T_3[6:0] ? myVec_24 : _GEN_10433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10435 = 7'h19 == _myNewVec_47_T_3[6:0] ? myVec_25 : _GEN_10434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10436 = 7'h1a == _myNewVec_47_T_3[6:0] ? myVec_26 : _GEN_10435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10437 = 7'h1b == _myNewVec_47_T_3[6:0] ? myVec_27 : _GEN_10436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10438 = 7'h1c == _myNewVec_47_T_3[6:0] ? myVec_28 : _GEN_10437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10439 = 7'h1d == _myNewVec_47_T_3[6:0] ? myVec_29 : _GEN_10438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10440 = 7'h1e == _myNewVec_47_T_3[6:0] ? myVec_30 : _GEN_10439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10441 = 7'h1f == _myNewVec_47_T_3[6:0] ? myVec_31 : _GEN_10440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10442 = 7'h20 == _myNewVec_47_T_3[6:0] ? myVec_32 : _GEN_10441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10443 = 7'h21 == _myNewVec_47_T_3[6:0] ? myVec_33 : _GEN_10442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10444 = 7'h22 == _myNewVec_47_T_3[6:0] ? myVec_34 : _GEN_10443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10445 = 7'h23 == _myNewVec_47_T_3[6:0] ? myVec_35 : _GEN_10444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10446 = 7'h24 == _myNewVec_47_T_3[6:0] ? myVec_36 : _GEN_10445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10447 = 7'h25 == _myNewVec_47_T_3[6:0] ? myVec_37 : _GEN_10446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10448 = 7'h26 == _myNewVec_47_T_3[6:0] ? myVec_38 : _GEN_10447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10449 = 7'h27 == _myNewVec_47_T_3[6:0] ? myVec_39 : _GEN_10448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10450 = 7'h28 == _myNewVec_47_T_3[6:0] ? myVec_40 : _GEN_10449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10451 = 7'h29 == _myNewVec_47_T_3[6:0] ? myVec_41 : _GEN_10450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10452 = 7'h2a == _myNewVec_47_T_3[6:0] ? myVec_42 : _GEN_10451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10453 = 7'h2b == _myNewVec_47_T_3[6:0] ? myVec_43 : _GEN_10452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10454 = 7'h2c == _myNewVec_47_T_3[6:0] ? myVec_44 : _GEN_10453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10455 = 7'h2d == _myNewVec_47_T_3[6:0] ? myVec_45 : _GEN_10454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10456 = 7'h2e == _myNewVec_47_T_3[6:0] ? myVec_46 : _GEN_10455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10457 = 7'h2f == _myNewVec_47_T_3[6:0] ? myVec_47 : _GEN_10456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10458 = 7'h30 == _myNewVec_47_T_3[6:0] ? myVec_48 : _GEN_10457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10459 = 7'h31 == _myNewVec_47_T_3[6:0] ? myVec_49 : _GEN_10458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10460 = 7'h32 == _myNewVec_47_T_3[6:0] ? myVec_50 : _GEN_10459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10461 = 7'h33 == _myNewVec_47_T_3[6:0] ? myVec_51 : _GEN_10460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10462 = 7'h34 == _myNewVec_47_T_3[6:0] ? myVec_52 : _GEN_10461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10463 = 7'h35 == _myNewVec_47_T_3[6:0] ? myVec_53 : _GEN_10462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10464 = 7'h36 == _myNewVec_47_T_3[6:0] ? myVec_54 : _GEN_10463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10465 = 7'h37 == _myNewVec_47_T_3[6:0] ? myVec_55 : _GEN_10464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10466 = 7'h38 == _myNewVec_47_T_3[6:0] ? myVec_56 : _GEN_10465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10467 = 7'h39 == _myNewVec_47_T_3[6:0] ? myVec_57 : _GEN_10466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10468 = 7'h3a == _myNewVec_47_T_3[6:0] ? myVec_58 : _GEN_10467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10469 = 7'h3b == _myNewVec_47_T_3[6:0] ? myVec_59 : _GEN_10468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10470 = 7'h3c == _myNewVec_47_T_3[6:0] ? myVec_60 : _GEN_10469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10471 = 7'h3d == _myNewVec_47_T_3[6:0] ? myVec_61 : _GEN_10470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10472 = 7'h3e == _myNewVec_47_T_3[6:0] ? myVec_62 : _GEN_10471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10473 = 7'h3f == _myNewVec_47_T_3[6:0] ? myVec_63 : _GEN_10472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10474 = 7'h40 == _myNewVec_47_T_3[6:0] ? myVec_64 : _GEN_10473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10475 = 7'h41 == _myNewVec_47_T_3[6:0] ? myVec_65 : _GEN_10474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10476 = 7'h42 == _myNewVec_47_T_3[6:0] ? myVec_66 : _GEN_10475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10477 = 7'h43 == _myNewVec_47_T_3[6:0] ? myVec_67 : _GEN_10476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10478 = 7'h44 == _myNewVec_47_T_3[6:0] ? myVec_68 : _GEN_10477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10479 = 7'h45 == _myNewVec_47_T_3[6:0] ? myVec_69 : _GEN_10478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10480 = 7'h46 == _myNewVec_47_T_3[6:0] ? myVec_70 : _GEN_10479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10481 = 7'h47 == _myNewVec_47_T_3[6:0] ? myVec_71 : _GEN_10480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10482 = 7'h48 == _myNewVec_47_T_3[6:0] ? myVec_72 : _GEN_10481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10483 = 7'h49 == _myNewVec_47_T_3[6:0] ? myVec_73 : _GEN_10482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10484 = 7'h4a == _myNewVec_47_T_3[6:0] ? myVec_74 : _GEN_10483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10485 = 7'h4b == _myNewVec_47_T_3[6:0] ? myVec_75 : _GEN_10484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10486 = 7'h4c == _myNewVec_47_T_3[6:0] ? myVec_76 : _GEN_10485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10487 = 7'h4d == _myNewVec_47_T_3[6:0] ? myVec_77 : _GEN_10486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10488 = 7'h4e == _myNewVec_47_T_3[6:0] ? myVec_78 : _GEN_10487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10489 = 7'h4f == _myNewVec_47_T_3[6:0] ? myVec_79 : _GEN_10488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10490 = 7'h50 == _myNewVec_47_T_3[6:0] ? myVec_80 : _GEN_10489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10491 = 7'h51 == _myNewVec_47_T_3[6:0] ? myVec_81 : _GEN_10490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10492 = 7'h52 == _myNewVec_47_T_3[6:0] ? myVec_82 : _GEN_10491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10493 = 7'h53 == _myNewVec_47_T_3[6:0] ? myVec_83 : _GEN_10492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10494 = 7'h54 == _myNewVec_47_T_3[6:0] ? myVec_84 : _GEN_10493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10495 = 7'h55 == _myNewVec_47_T_3[6:0] ? myVec_85 : _GEN_10494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10496 = 7'h56 == _myNewVec_47_T_3[6:0] ? myVec_86 : _GEN_10495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10497 = 7'h57 == _myNewVec_47_T_3[6:0] ? myVec_87 : _GEN_10496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10498 = 7'h58 == _myNewVec_47_T_3[6:0] ? myVec_88 : _GEN_10497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10499 = 7'h59 == _myNewVec_47_T_3[6:0] ? myVec_89 : _GEN_10498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10500 = 7'h5a == _myNewVec_47_T_3[6:0] ? myVec_90 : _GEN_10499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10501 = 7'h5b == _myNewVec_47_T_3[6:0] ? myVec_91 : _GEN_10500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10502 = 7'h5c == _myNewVec_47_T_3[6:0] ? myVec_92 : _GEN_10501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10503 = 7'h5d == _myNewVec_47_T_3[6:0] ? myVec_93 : _GEN_10502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10504 = 7'h5e == _myNewVec_47_T_3[6:0] ? myVec_94 : _GEN_10503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10505 = 7'h5f == _myNewVec_47_T_3[6:0] ? myVec_95 : _GEN_10504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10506 = 7'h60 == _myNewVec_47_T_3[6:0] ? myVec_96 : _GEN_10505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10507 = 7'h61 == _myNewVec_47_T_3[6:0] ? myVec_97 : _GEN_10506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10508 = 7'h62 == _myNewVec_47_T_3[6:0] ? myVec_98 : _GEN_10507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10509 = 7'h63 == _myNewVec_47_T_3[6:0] ? myVec_99 : _GEN_10508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10510 = 7'h64 == _myNewVec_47_T_3[6:0] ? myVec_100 : _GEN_10509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10511 = 7'h65 == _myNewVec_47_T_3[6:0] ? myVec_101 : _GEN_10510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10512 = 7'h66 == _myNewVec_47_T_3[6:0] ? myVec_102 : _GEN_10511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10513 = 7'h67 == _myNewVec_47_T_3[6:0] ? myVec_103 : _GEN_10512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10514 = 7'h68 == _myNewVec_47_T_3[6:0] ? myVec_104 : _GEN_10513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10515 = 7'h69 == _myNewVec_47_T_3[6:0] ? myVec_105 : _GEN_10514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10516 = 7'h6a == _myNewVec_47_T_3[6:0] ? myVec_106 : _GEN_10515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10517 = 7'h6b == _myNewVec_47_T_3[6:0] ? myVec_107 : _GEN_10516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10518 = 7'h6c == _myNewVec_47_T_3[6:0] ? myVec_108 : _GEN_10517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10519 = 7'h6d == _myNewVec_47_T_3[6:0] ? myVec_109 : _GEN_10518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10520 = 7'h6e == _myNewVec_47_T_3[6:0] ? myVec_110 : _GEN_10519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10521 = 7'h6f == _myNewVec_47_T_3[6:0] ? myVec_111 : _GEN_10520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10522 = 7'h70 == _myNewVec_47_T_3[6:0] ? myVec_112 : _GEN_10521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10523 = 7'h71 == _myNewVec_47_T_3[6:0] ? myVec_113 : _GEN_10522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10524 = 7'h72 == _myNewVec_47_T_3[6:0] ? myVec_114 : _GEN_10523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10525 = 7'h73 == _myNewVec_47_T_3[6:0] ? myVec_115 : _GEN_10524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10526 = 7'h74 == _myNewVec_47_T_3[6:0] ? myVec_116 : _GEN_10525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10527 = 7'h75 == _myNewVec_47_T_3[6:0] ? myVec_117 : _GEN_10526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10528 = 7'h76 == _myNewVec_47_T_3[6:0] ? myVec_118 : _GEN_10527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10529 = 7'h77 == _myNewVec_47_T_3[6:0] ? myVec_119 : _GEN_10528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10530 = 7'h78 == _myNewVec_47_T_3[6:0] ? myVec_120 : _GEN_10529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10531 = 7'h79 == _myNewVec_47_T_3[6:0] ? myVec_121 : _GEN_10530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10532 = 7'h7a == _myNewVec_47_T_3[6:0] ? myVec_122 : _GEN_10531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10533 = 7'h7b == _myNewVec_47_T_3[6:0] ? myVec_123 : _GEN_10532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10534 = 7'h7c == _myNewVec_47_T_3[6:0] ? myVec_124 : _GEN_10533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10535 = 7'h7d == _myNewVec_47_T_3[6:0] ? myVec_125 : _GEN_10534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10536 = 7'h7e == _myNewVec_47_T_3[6:0] ? myVec_126 : _GEN_10535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_47 = 7'h7f == _myNewVec_47_T_3[6:0] ? myVec_127 : _GEN_10536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_46_T_3 = _myNewVec_127_T_1 + 16'h51; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_10539 = 7'h1 == _myNewVec_46_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10540 = 7'h2 == _myNewVec_46_T_3[6:0] ? myVec_2 : _GEN_10539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10541 = 7'h3 == _myNewVec_46_T_3[6:0] ? myVec_3 : _GEN_10540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10542 = 7'h4 == _myNewVec_46_T_3[6:0] ? myVec_4 : _GEN_10541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10543 = 7'h5 == _myNewVec_46_T_3[6:0] ? myVec_5 : _GEN_10542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10544 = 7'h6 == _myNewVec_46_T_3[6:0] ? myVec_6 : _GEN_10543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10545 = 7'h7 == _myNewVec_46_T_3[6:0] ? myVec_7 : _GEN_10544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10546 = 7'h8 == _myNewVec_46_T_3[6:0] ? myVec_8 : _GEN_10545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10547 = 7'h9 == _myNewVec_46_T_3[6:0] ? myVec_9 : _GEN_10546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10548 = 7'ha == _myNewVec_46_T_3[6:0] ? myVec_10 : _GEN_10547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10549 = 7'hb == _myNewVec_46_T_3[6:0] ? myVec_11 : _GEN_10548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10550 = 7'hc == _myNewVec_46_T_3[6:0] ? myVec_12 : _GEN_10549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10551 = 7'hd == _myNewVec_46_T_3[6:0] ? myVec_13 : _GEN_10550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10552 = 7'he == _myNewVec_46_T_3[6:0] ? myVec_14 : _GEN_10551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10553 = 7'hf == _myNewVec_46_T_3[6:0] ? myVec_15 : _GEN_10552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10554 = 7'h10 == _myNewVec_46_T_3[6:0] ? myVec_16 : _GEN_10553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10555 = 7'h11 == _myNewVec_46_T_3[6:0] ? myVec_17 : _GEN_10554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10556 = 7'h12 == _myNewVec_46_T_3[6:0] ? myVec_18 : _GEN_10555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10557 = 7'h13 == _myNewVec_46_T_3[6:0] ? myVec_19 : _GEN_10556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10558 = 7'h14 == _myNewVec_46_T_3[6:0] ? myVec_20 : _GEN_10557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10559 = 7'h15 == _myNewVec_46_T_3[6:0] ? myVec_21 : _GEN_10558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10560 = 7'h16 == _myNewVec_46_T_3[6:0] ? myVec_22 : _GEN_10559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10561 = 7'h17 == _myNewVec_46_T_3[6:0] ? myVec_23 : _GEN_10560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10562 = 7'h18 == _myNewVec_46_T_3[6:0] ? myVec_24 : _GEN_10561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10563 = 7'h19 == _myNewVec_46_T_3[6:0] ? myVec_25 : _GEN_10562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10564 = 7'h1a == _myNewVec_46_T_3[6:0] ? myVec_26 : _GEN_10563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10565 = 7'h1b == _myNewVec_46_T_3[6:0] ? myVec_27 : _GEN_10564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10566 = 7'h1c == _myNewVec_46_T_3[6:0] ? myVec_28 : _GEN_10565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10567 = 7'h1d == _myNewVec_46_T_3[6:0] ? myVec_29 : _GEN_10566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10568 = 7'h1e == _myNewVec_46_T_3[6:0] ? myVec_30 : _GEN_10567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10569 = 7'h1f == _myNewVec_46_T_3[6:0] ? myVec_31 : _GEN_10568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10570 = 7'h20 == _myNewVec_46_T_3[6:0] ? myVec_32 : _GEN_10569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10571 = 7'h21 == _myNewVec_46_T_3[6:0] ? myVec_33 : _GEN_10570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10572 = 7'h22 == _myNewVec_46_T_3[6:0] ? myVec_34 : _GEN_10571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10573 = 7'h23 == _myNewVec_46_T_3[6:0] ? myVec_35 : _GEN_10572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10574 = 7'h24 == _myNewVec_46_T_3[6:0] ? myVec_36 : _GEN_10573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10575 = 7'h25 == _myNewVec_46_T_3[6:0] ? myVec_37 : _GEN_10574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10576 = 7'h26 == _myNewVec_46_T_3[6:0] ? myVec_38 : _GEN_10575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10577 = 7'h27 == _myNewVec_46_T_3[6:0] ? myVec_39 : _GEN_10576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10578 = 7'h28 == _myNewVec_46_T_3[6:0] ? myVec_40 : _GEN_10577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10579 = 7'h29 == _myNewVec_46_T_3[6:0] ? myVec_41 : _GEN_10578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10580 = 7'h2a == _myNewVec_46_T_3[6:0] ? myVec_42 : _GEN_10579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10581 = 7'h2b == _myNewVec_46_T_3[6:0] ? myVec_43 : _GEN_10580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10582 = 7'h2c == _myNewVec_46_T_3[6:0] ? myVec_44 : _GEN_10581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10583 = 7'h2d == _myNewVec_46_T_3[6:0] ? myVec_45 : _GEN_10582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10584 = 7'h2e == _myNewVec_46_T_3[6:0] ? myVec_46 : _GEN_10583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10585 = 7'h2f == _myNewVec_46_T_3[6:0] ? myVec_47 : _GEN_10584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10586 = 7'h30 == _myNewVec_46_T_3[6:0] ? myVec_48 : _GEN_10585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10587 = 7'h31 == _myNewVec_46_T_3[6:0] ? myVec_49 : _GEN_10586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10588 = 7'h32 == _myNewVec_46_T_3[6:0] ? myVec_50 : _GEN_10587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10589 = 7'h33 == _myNewVec_46_T_3[6:0] ? myVec_51 : _GEN_10588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10590 = 7'h34 == _myNewVec_46_T_3[6:0] ? myVec_52 : _GEN_10589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10591 = 7'h35 == _myNewVec_46_T_3[6:0] ? myVec_53 : _GEN_10590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10592 = 7'h36 == _myNewVec_46_T_3[6:0] ? myVec_54 : _GEN_10591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10593 = 7'h37 == _myNewVec_46_T_3[6:0] ? myVec_55 : _GEN_10592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10594 = 7'h38 == _myNewVec_46_T_3[6:0] ? myVec_56 : _GEN_10593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10595 = 7'h39 == _myNewVec_46_T_3[6:0] ? myVec_57 : _GEN_10594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10596 = 7'h3a == _myNewVec_46_T_3[6:0] ? myVec_58 : _GEN_10595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10597 = 7'h3b == _myNewVec_46_T_3[6:0] ? myVec_59 : _GEN_10596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10598 = 7'h3c == _myNewVec_46_T_3[6:0] ? myVec_60 : _GEN_10597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10599 = 7'h3d == _myNewVec_46_T_3[6:0] ? myVec_61 : _GEN_10598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10600 = 7'h3e == _myNewVec_46_T_3[6:0] ? myVec_62 : _GEN_10599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10601 = 7'h3f == _myNewVec_46_T_3[6:0] ? myVec_63 : _GEN_10600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10602 = 7'h40 == _myNewVec_46_T_3[6:0] ? myVec_64 : _GEN_10601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10603 = 7'h41 == _myNewVec_46_T_3[6:0] ? myVec_65 : _GEN_10602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10604 = 7'h42 == _myNewVec_46_T_3[6:0] ? myVec_66 : _GEN_10603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10605 = 7'h43 == _myNewVec_46_T_3[6:0] ? myVec_67 : _GEN_10604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10606 = 7'h44 == _myNewVec_46_T_3[6:0] ? myVec_68 : _GEN_10605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10607 = 7'h45 == _myNewVec_46_T_3[6:0] ? myVec_69 : _GEN_10606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10608 = 7'h46 == _myNewVec_46_T_3[6:0] ? myVec_70 : _GEN_10607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10609 = 7'h47 == _myNewVec_46_T_3[6:0] ? myVec_71 : _GEN_10608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10610 = 7'h48 == _myNewVec_46_T_3[6:0] ? myVec_72 : _GEN_10609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10611 = 7'h49 == _myNewVec_46_T_3[6:0] ? myVec_73 : _GEN_10610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10612 = 7'h4a == _myNewVec_46_T_3[6:0] ? myVec_74 : _GEN_10611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10613 = 7'h4b == _myNewVec_46_T_3[6:0] ? myVec_75 : _GEN_10612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10614 = 7'h4c == _myNewVec_46_T_3[6:0] ? myVec_76 : _GEN_10613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10615 = 7'h4d == _myNewVec_46_T_3[6:0] ? myVec_77 : _GEN_10614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10616 = 7'h4e == _myNewVec_46_T_3[6:0] ? myVec_78 : _GEN_10615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10617 = 7'h4f == _myNewVec_46_T_3[6:0] ? myVec_79 : _GEN_10616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10618 = 7'h50 == _myNewVec_46_T_3[6:0] ? myVec_80 : _GEN_10617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10619 = 7'h51 == _myNewVec_46_T_3[6:0] ? myVec_81 : _GEN_10618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10620 = 7'h52 == _myNewVec_46_T_3[6:0] ? myVec_82 : _GEN_10619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10621 = 7'h53 == _myNewVec_46_T_3[6:0] ? myVec_83 : _GEN_10620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10622 = 7'h54 == _myNewVec_46_T_3[6:0] ? myVec_84 : _GEN_10621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10623 = 7'h55 == _myNewVec_46_T_3[6:0] ? myVec_85 : _GEN_10622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10624 = 7'h56 == _myNewVec_46_T_3[6:0] ? myVec_86 : _GEN_10623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10625 = 7'h57 == _myNewVec_46_T_3[6:0] ? myVec_87 : _GEN_10624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10626 = 7'h58 == _myNewVec_46_T_3[6:0] ? myVec_88 : _GEN_10625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10627 = 7'h59 == _myNewVec_46_T_3[6:0] ? myVec_89 : _GEN_10626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10628 = 7'h5a == _myNewVec_46_T_3[6:0] ? myVec_90 : _GEN_10627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10629 = 7'h5b == _myNewVec_46_T_3[6:0] ? myVec_91 : _GEN_10628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10630 = 7'h5c == _myNewVec_46_T_3[6:0] ? myVec_92 : _GEN_10629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10631 = 7'h5d == _myNewVec_46_T_3[6:0] ? myVec_93 : _GEN_10630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10632 = 7'h5e == _myNewVec_46_T_3[6:0] ? myVec_94 : _GEN_10631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10633 = 7'h5f == _myNewVec_46_T_3[6:0] ? myVec_95 : _GEN_10632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10634 = 7'h60 == _myNewVec_46_T_3[6:0] ? myVec_96 : _GEN_10633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10635 = 7'h61 == _myNewVec_46_T_3[6:0] ? myVec_97 : _GEN_10634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10636 = 7'h62 == _myNewVec_46_T_3[6:0] ? myVec_98 : _GEN_10635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10637 = 7'h63 == _myNewVec_46_T_3[6:0] ? myVec_99 : _GEN_10636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10638 = 7'h64 == _myNewVec_46_T_3[6:0] ? myVec_100 : _GEN_10637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10639 = 7'h65 == _myNewVec_46_T_3[6:0] ? myVec_101 : _GEN_10638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10640 = 7'h66 == _myNewVec_46_T_3[6:0] ? myVec_102 : _GEN_10639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10641 = 7'h67 == _myNewVec_46_T_3[6:0] ? myVec_103 : _GEN_10640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10642 = 7'h68 == _myNewVec_46_T_3[6:0] ? myVec_104 : _GEN_10641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10643 = 7'h69 == _myNewVec_46_T_3[6:0] ? myVec_105 : _GEN_10642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10644 = 7'h6a == _myNewVec_46_T_3[6:0] ? myVec_106 : _GEN_10643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10645 = 7'h6b == _myNewVec_46_T_3[6:0] ? myVec_107 : _GEN_10644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10646 = 7'h6c == _myNewVec_46_T_3[6:0] ? myVec_108 : _GEN_10645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10647 = 7'h6d == _myNewVec_46_T_3[6:0] ? myVec_109 : _GEN_10646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10648 = 7'h6e == _myNewVec_46_T_3[6:0] ? myVec_110 : _GEN_10647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10649 = 7'h6f == _myNewVec_46_T_3[6:0] ? myVec_111 : _GEN_10648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10650 = 7'h70 == _myNewVec_46_T_3[6:0] ? myVec_112 : _GEN_10649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10651 = 7'h71 == _myNewVec_46_T_3[6:0] ? myVec_113 : _GEN_10650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10652 = 7'h72 == _myNewVec_46_T_3[6:0] ? myVec_114 : _GEN_10651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10653 = 7'h73 == _myNewVec_46_T_3[6:0] ? myVec_115 : _GEN_10652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10654 = 7'h74 == _myNewVec_46_T_3[6:0] ? myVec_116 : _GEN_10653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10655 = 7'h75 == _myNewVec_46_T_3[6:0] ? myVec_117 : _GEN_10654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10656 = 7'h76 == _myNewVec_46_T_3[6:0] ? myVec_118 : _GEN_10655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10657 = 7'h77 == _myNewVec_46_T_3[6:0] ? myVec_119 : _GEN_10656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10658 = 7'h78 == _myNewVec_46_T_3[6:0] ? myVec_120 : _GEN_10657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10659 = 7'h79 == _myNewVec_46_T_3[6:0] ? myVec_121 : _GEN_10658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10660 = 7'h7a == _myNewVec_46_T_3[6:0] ? myVec_122 : _GEN_10659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10661 = 7'h7b == _myNewVec_46_T_3[6:0] ? myVec_123 : _GEN_10660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10662 = 7'h7c == _myNewVec_46_T_3[6:0] ? myVec_124 : _GEN_10661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10663 = 7'h7d == _myNewVec_46_T_3[6:0] ? myVec_125 : _GEN_10662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10664 = 7'h7e == _myNewVec_46_T_3[6:0] ? myVec_126 : _GEN_10663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_46 = 7'h7f == _myNewVec_46_T_3[6:0] ? myVec_127 : _GEN_10664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_45_T_3 = _myNewVec_127_T_1 + 16'h52; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_10667 = 7'h1 == _myNewVec_45_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10668 = 7'h2 == _myNewVec_45_T_3[6:0] ? myVec_2 : _GEN_10667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10669 = 7'h3 == _myNewVec_45_T_3[6:0] ? myVec_3 : _GEN_10668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10670 = 7'h4 == _myNewVec_45_T_3[6:0] ? myVec_4 : _GEN_10669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10671 = 7'h5 == _myNewVec_45_T_3[6:0] ? myVec_5 : _GEN_10670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10672 = 7'h6 == _myNewVec_45_T_3[6:0] ? myVec_6 : _GEN_10671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10673 = 7'h7 == _myNewVec_45_T_3[6:0] ? myVec_7 : _GEN_10672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10674 = 7'h8 == _myNewVec_45_T_3[6:0] ? myVec_8 : _GEN_10673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10675 = 7'h9 == _myNewVec_45_T_3[6:0] ? myVec_9 : _GEN_10674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10676 = 7'ha == _myNewVec_45_T_3[6:0] ? myVec_10 : _GEN_10675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10677 = 7'hb == _myNewVec_45_T_3[6:0] ? myVec_11 : _GEN_10676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10678 = 7'hc == _myNewVec_45_T_3[6:0] ? myVec_12 : _GEN_10677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10679 = 7'hd == _myNewVec_45_T_3[6:0] ? myVec_13 : _GEN_10678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10680 = 7'he == _myNewVec_45_T_3[6:0] ? myVec_14 : _GEN_10679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10681 = 7'hf == _myNewVec_45_T_3[6:0] ? myVec_15 : _GEN_10680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10682 = 7'h10 == _myNewVec_45_T_3[6:0] ? myVec_16 : _GEN_10681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10683 = 7'h11 == _myNewVec_45_T_3[6:0] ? myVec_17 : _GEN_10682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10684 = 7'h12 == _myNewVec_45_T_3[6:0] ? myVec_18 : _GEN_10683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10685 = 7'h13 == _myNewVec_45_T_3[6:0] ? myVec_19 : _GEN_10684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10686 = 7'h14 == _myNewVec_45_T_3[6:0] ? myVec_20 : _GEN_10685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10687 = 7'h15 == _myNewVec_45_T_3[6:0] ? myVec_21 : _GEN_10686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10688 = 7'h16 == _myNewVec_45_T_3[6:0] ? myVec_22 : _GEN_10687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10689 = 7'h17 == _myNewVec_45_T_3[6:0] ? myVec_23 : _GEN_10688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10690 = 7'h18 == _myNewVec_45_T_3[6:0] ? myVec_24 : _GEN_10689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10691 = 7'h19 == _myNewVec_45_T_3[6:0] ? myVec_25 : _GEN_10690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10692 = 7'h1a == _myNewVec_45_T_3[6:0] ? myVec_26 : _GEN_10691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10693 = 7'h1b == _myNewVec_45_T_3[6:0] ? myVec_27 : _GEN_10692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10694 = 7'h1c == _myNewVec_45_T_3[6:0] ? myVec_28 : _GEN_10693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10695 = 7'h1d == _myNewVec_45_T_3[6:0] ? myVec_29 : _GEN_10694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10696 = 7'h1e == _myNewVec_45_T_3[6:0] ? myVec_30 : _GEN_10695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10697 = 7'h1f == _myNewVec_45_T_3[6:0] ? myVec_31 : _GEN_10696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10698 = 7'h20 == _myNewVec_45_T_3[6:0] ? myVec_32 : _GEN_10697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10699 = 7'h21 == _myNewVec_45_T_3[6:0] ? myVec_33 : _GEN_10698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10700 = 7'h22 == _myNewVec_45_T_3[6:0] ? myVec_34 : _GEN_10699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10701 = 7'h23 == _myNewVec_45_T_3[6:0] ? myVec_35 : _GEN_10700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10702 = 7'h24 == _myNewVec_45_T_3[6:0] ? myVec_36 : _GEN_10701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10703 = 7'h25 == _myNewVec_45_T_3[6:0] ? myVec_37 : _GEN_10702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10704 = 7'h26 == _myNewVec_45_T_3[6:0] ? myVec_38 : _GEN_10703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10705 = 7'h27 == _myNewVec_45_T_3[6:0] ? myVec_39 : _GEN_10704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10706 = 7'h28 == _myNewVec_45_T_3[6:0] ? myVec_40 : _GEN_10705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10707 = 7'h29 == _myNewVec_45_T_3[6:0] ? myVec_41 : _GEN_10706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10708 = 7'h2a == _myNewVec_45_T_3[6:0] ? myVec_42 : _GEN_10707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10709 = 7'h2b == _myNewVec_45_T_3[6:0] ? myVec_43 : _GEN_10708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10710 = 7'h2c == _myNewVec_45_T_3[6:0] ? myVec_44 : _GEN_10709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10711 = 7'h2d == _myNewVec_45_T_3[6:0] ? myVec_45 : _GEN_10710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10712 = 7'h2e == _myNewVec_45_T_3[6:0] ? myVec_46 : _GEN_10711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10713 = 7'h2f == _myNewVec_45_T_3[6:0] ? myVec_47 : _GEN_10712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10714 = 7'h30 == _myNewVec_45_T_3[6:0] ? myVec_48 : _GEN_10713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10715 = 7'h31 == _myNewVec_45_T_3[6:0] ? myVec_49 : _GEN_10714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10716 = 7'h32 == _myNewVec_45_T_3[6:0] ? myVec_50 : _GEN_10715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10717 = 7'h33 == _myNewVec_45_T_3[6:0] ? myVec_51 : _GEN_10716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10718 = 7'h34 == _myNewVec_45_T_3[6:0] ? myVec_52 : _GEN_10717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10719 = 7'h35 == _myNewVec_45_T_3[6:0] ? myVec_53 : _GEN_10718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10720 = 7'h36 == _myNewVec_45_T_3[6:0] ? myVec_54 : _GEN_10719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10721 = 7'h37 == _myNewVec_45_T_3[6:0] ? myVec_55 : _GEN_10720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10722 = 7'h38 == _myNewVec_45_T_3[6:0] ? myVec_56 : _GEN_10721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10723 = 7'h39 == _myNewVec_45_T_3[6:0] ? myVec_57 : _GEN_10722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10724 = 7'h3a == _myNewVec_45_T_3[6:0] ? myVec_58 : _GEN_10723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10725 = 7'h3b == _myNewVec_45_T_3[6:0] ? myVec_59 : _GEN_10724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10726 = 7'h3c == _myNewVec_45_T_3[6:0] ? myVec_60 : _GEN_10725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10727 = 7'h3d == _myNewVec_45_T_3[6:0] ? myVec_61 : _GEN_10726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10728 = 7'h3e == _myNewVec_45_T_3[6:0] ? myVec_62 : _GEN_10727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10729 = 7'h3f == _myNewVec_45_T_3[6:0] ? myVec_63 : _GEN_10728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10730 = 7'h40 == _myNewVec_45_T_3[6:0] ? myVec_64 : _GEN_10729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10731 = 7'h41 == _myNewVec_45_T_3[6:0] ? myVec_65 : _GEN_10730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10732 = 7'h42 == _myNewVec_45_T_3[6:0] ? myVec_66 : _GEN_10731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10733 = 7'h43 == _myNewVec_45_T_3[6:0] ? myVec_67 : _GEN_10732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10734 = 7'h44 == _myNewVec_45_T_3[6:0] ? myVec_68 : _GEN_10733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10735 = 7'h45 == _myNewVec_45_T_3[6:0] ? myVec_69 : _GEN_10734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10736 = 7'h46 == _myNewVec_45_T_3[6:0] ? myVec_70 : _GEN_10735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10737 = 7'h47 == _myNewVec_45_T_3[6:0] ? myVec_71 : _GEN_10736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10738 = 7'h48 == _myNewVec_45_T_3[6:0] ? myVec_72 : _GEN_10737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10739 = 7'h49 == _myNewVec_45_T_3[6:0] ? myVec_73 : _GEN_10738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10740 = 7'h4a == _myNewVec_45_T_3[6:0] ? myVec_74 : _GEN_10739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10741 = 7'h4b == _myNewVec_45_T_3[6:0] ? myVec_75 : _GEN_10740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10742 = 7'h4c == _myNewVec_45_T_3[6:0] ? myVec_76 : _GEN_10741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10743 = 7'h4d == _myNewVec_45_T_3[6:0] ? myVec_77 : _GEN_10742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10744 = 7'h4e == _myNewVec_45_T_3[6:0] ? myVec_78 : _GEN_10743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10745 = 7'h4f == _myNewVec_45_T_3[6:0] ? myVec_79 : _GEN_10744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10746 = 7'h50 == _myNewVec_45_T_3[6:0] ? myVec_80 : _GEN_10745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10747 = 7'h51 == _myNewVec_45_T_3[6:0] ? myVec_81 : _GEN_10746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10748 = 7'h52 == _myNewVec_45_T_3[6:0] ? myVec_82 : _GEN_10747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10749 = 7'h53 == _myNewVec_45_T_3[6:0] ? myVec_83 : _GEN_10748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10750 = 7'h54 == _myNewVec_45_T_3[6:0] ? myVec_84 : _GEN_10749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10751 = 7'h55 == _myNewVec_45_T_3[6:0] ? myVec_85 : _GEN_10750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10752 = 7'h56 == _myNewVec_45_T_3[6:0] ? myVec_86 : _GEN_10751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10753 = 7'h57 == _myNewVec_45_T_3[6:0] ? myVec_87 : _GEN_10752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10754 = 7'h58 == _myNewVec_45_T_3[6:0] ? myVec_88 : _GEN_10753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10755 = 7'h59 == _myNewVec_45_T_3[6:0] ? myVec_89 : _GEN_10754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10756 = 7'h5a == _myNewVec_45_T_3[6:0] ? myVec_90 : _GEN_10755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10757 = 7'h5b == _myNewVec_45_T_3[6:0] ? myVec_91 : _GEN_10756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10758 = 7'h5c == _myNewVec_45_T_3[6:0] ? myVec_92 : _GEN_10757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10759 = 7'h5d == _myNewVec_45_T_3[6:0] ? myVec_93 : _GEN_10758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10760 = 7'h5e == _myNewVec_45_T_3[6:0] ? myVec_94 : _GEN_10759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10761 = 7'h5f == _myNewVec_45_T_3[6:0] ? myVec_95 : _GEN_10760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10762 = 7'h60 == _myNewVec_45_T_3[6:0] ? myVec_96 : _GEN_10761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10763 = 7'h61 == _myNewVec_45_T_3[6:0] ? myVec_97 : _GEN_10762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10764 = 7'h62 == _myNewVec_45_T_3[6:0] ? myVec_98 : _GEN_10763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10765 = 7'h63 == _myNewVec_45_T_3[6:0] ? myVec_99 : _GEN_10764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10766 = 7'h64 == _myNewVec_45_T_3[6:0] ? myVec_100 : _GEN_10765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10767 = 7'h65 == _myNewVec_45_T_3[6:0] ? myVec_101 : _GEN_10766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10768 = 7'h66 == _myNewVec_45_T_3[6:0] ? myVec_102 : _GEN_10767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10769 = 7'h67 == _myNewVec_45_T_3[6:0] ? myVec_103 : _GEN_10768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10770 = 7'h68 == _myNewVec_45_T_3[6:0] ? myVec_104 : _GEN_10769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10771 = 7'h69 == _myNewVec_45_T_3[6:0] ? myVec_105 : _GEN_10770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10772 = 7'h6a == _myNewVec_45_T_3[6:0] ? myVec_106 : _GEN_10771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10773 = 7'h6b == _myNewVec_45_T_3[6:0] ? myVec_107 : _GEN_10772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10774 = 7'h6c == _myNewVec_45_T_3[6:0] ? myVec_108 : _GEN_10773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10775 = 7'h6d == _myNewVec_45_T_3[6:0] ? myVec_109 : _GEN_10774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10776 = 7'h6e == _myNewVec_45_T_3[6:0] ? myVec_110 : _GEN_10775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10777 = 7'h6f == _myNewVec_45_T_3[6:0] ? myVec_111 : _GEN_10776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10778 = 7'h70 == _myNewVec_45_T_3[6:0] ? myVec_112 : _GEN_10777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10779 = 7'h71 == _myNewVec_45_T_3[6:0] ? myVec_113 : _GEN_10778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10780 = 7'h72 == _myNewVec_45_T_3[6:0] ? myVec_114 : _GEN_10779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10781 = 7'h73 == _myNewVec_45_T_3[6:0] ? myVec_115 : _GEN_10780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10782 = 7'h74 == _myNewVec_45_T_3[6:0] ? myVec_116 : _GEN_10781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10783 = 7'h75 == _myNewVec_45_T_3[6:0] ? myVec_117 : _GEN_10782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10784 = 7'h76 == _myNewVec_45_T_3[6:0] ? myVec_118 : _GEN_10783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10785 = 7'h77 == _myNewVec_45_T_3[6:0] ? myVec_119 : _GEN_10784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10786 = 7'h78 == _myNewVec_45_T_3[6:0] ? myVec_120 : _GEN_10785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10787 = 7'h79 == _myNewVec_45_T_3[6:0] ? myVec_121 : _GEN_10786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10788 = 7'h7a == _myNewVec_45_T_3[6:0] ? myVec_122 : _GEN_10787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10789 = 7'h7b == _myNewVec_45_T_3[6:0] ? myVec_123 : _GEN_10788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10790 = 7'h7c == _myNewVec_45_T_3[6:0] ? myVec_124 : _GEN_10789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10791 = 7'h7d == _myNewVec_45_T_3[6:0] ? myVec_125 : _GEN_10790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10792 = 7'h7e == _myNewVec_45_T_3[6:0] ? myVec_126 : _GEN_10791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_45 = 7'h7f == _myNewVec_45_T_3[6:0] ? myVec_127 : _GEN_10792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_44_T_3 = _myNewVec_127_T_1 + 16'h53; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_10795 = 7'h1 == _myNewVec_44_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10796 = 7'h2 == _myNewVec_44_T_3[6:0] ? myVec_2 : _GEN_10795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10797 = 7'h3 == _myNewVec_44_T_3[6:0] ? myVec_3 : _GEN_10796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10798 = 7'h4 == _myNewVec_44_T_3[6:0] ? myVec_4 : _GEN_10797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10799 = 7'h5 == _myNewVec_44_T_3[6:0] ? myVec_5 : _GEN_10798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10800 = 7'h6 == _myNewVec_44_T_3[6:0] ? myVec_6 : _GEN_10799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10801 = 7'h7 == _myNewVec_44_T_3[6:0] ? myVec_7 : _GEN_10800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10802 = 7'h8 == _myNewVec_44_T_3[6:0] ? myVec_8 : _GEN_10801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10803 = 7'h9 == _myNewVec_44_T_3[6:0] ? myVec_9 : _GEN_10802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10804 = 7'ha == _myNewVec_44_T_3[6:0] ? myVec_10 : _GEN_10803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10805 = 7'hb == _myNewVec_44_T_3[6:0] ? myVec_11 : _GEN_10804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10806 = 7'hc == _myNewVec_44_T_3[6:0] ? myVec_12 : _GEN_10805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10807 = 7'hd == _myNewVec_44_T_3[6:0] ? myVec_13 : _GEN_10806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10808 = 7'he == _myNewVec_44_T_3[6:0] ? myVec_14 : _GEN_10807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10809 = 7'hf == _myNewVec_44_T_3[6:0] ? myVec_15 : _GEN_10808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10810 = 7'h10 == _myNewVec_44_T_3[6:0] ? myVec_16 : _GEN_10809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10811 = 7'h11 == _myNewVec_44_T_3[6:0] ? myVec_17 : _GEN_10810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10812 = 7'h12 == _myNewVec_44_T_3[6:0] ? myVec_18 : _GEN_10811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10813 = 7'h13 == _myNewVec_44_T_3[6:0] ? myVec_19 : _GEN_10812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10814 = 7'h14 == _myNewVec_44_T_3[6:0] ? myVec_20 : _GEN_10813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10815 = 7'h15 == _myNewVec_44_T_3[6:0] ? myVec_21 : _GEN_10814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10816 = 7'h16 == _myNewVec_44_T_3[6:0] ? myVec_22 : _GEN_10815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10817 = 7'h17 == _myNewVec_44_T_3[6:0] ? myVec_23 : _GEN_10816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10818 = 7'h18 == _myNewVec_44_T_3[6:0] ? myVec_24 : _GEN_10817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10819 = 7'h19 == _myNewVec_44_T_3[6:0] ? myVec_25 : _GEN_10818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10820 = 7'h1a == _myNewVec_44_T_3[6:0] ? myVec_26 : _GEN_10819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10821 = 7'h1b == _myNewVec_44_T_3[6:0] ? myVec_27 : _GEN_10820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10822 = 7'h1c == _myNewVec_44_T_3[6:0] ? myVec_28 : _GEN_10821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10823 = 7'h1d == _myNewVec_44_T_3[6:0] ? myVec_29 : _GEN_10822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10824 = 7'h1e == _myNewVec_44_T_3[6:0] ? myVec_30 : _GEN_10823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10825 = 7'h1f == _myNewVec_44_T_3[6:0] ? myVec_31 : _GEN_10824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10826 = 7'h20 == _myNewVec_44_T_3[6:0] ? myVec_32 : _GEN_10825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10827 = 7'h21 == _myNewVec_44_T_3[6:0] ? myVec_33 : _GEN_10826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10828 = 7'h22 == _myNewVec_44_T_3[6:0] ? myVec_34 : _GEN_10827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10829 = 7'h23 == _myNewVec_44_T_3[6:0] ? myVec_35 : _GEN_10828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10830 = 7'h24 == _myNewVec_44_T_3[6:0] ? myVec_36 : _GEN_10829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10831 = 7'h25 == _myNewVec_44_T_3[6:0] ? myVec_37 : _GEN_10830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10832 = 7'h26 == _myNewVec_44_T_3[6:0] ? myVec_38 : _GEN_10831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10833 = 7'h27 == _myNewVec_44_T_3[6:0] ? myVec_39 : _GEN_10832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10834 = 7'h28 == _myNewVec_44_T_3[6:0] ? myVec_40 : _GEN_10833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10835 = 7'h29 == _myNewVec_44_T_3[6:0] ? myVec_41 : _GEN_10834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10836 = 7'h2a == _myNewVec_44_T_3[6:0] ? myVec_42 : _GEN_10835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10837 = 7'h2b == _myNewVec_44_T_3[6:0] ? myVec_43 : _GEN_10836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10838 = 7'h2c == _myNewVec_44_T_3[6:0] ? myVec_44 : _GEN_10837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10839 = 7'h2d == _myNewVec_44_T_3[6:0] ? myVec_45 : _GEN_10838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10840 = 7'h2e == _myNewVec_44_T_3[6:0] ? myVec_46 : _GEN_10839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10841 = 7'h2f == _myNewVec_44_T_3[6:0] ? myVec_47 : _GEN_10840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10842 = 7'h30 == _myNewVec_44_T_3[6:0] ? myVec_48 : _GEN_10841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10843 = 7'h31 == _myNewVec_44_T_3[6:0] ? myVec_49 : _GEN_10842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10844 = 7'h32 == _myNewVec_44_T_3[6:0] ? myVec_50 : _GEN_10843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10845 = 7'h33 == _myNewVec_44_T_3[6:0] ? myVec_51 : _GEN_10844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10846 = 7'h34 == _myNewVec_44_T_3[6:0] ? myVec_52 : _GEN_10845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10847 = 7'h35 == _myNewVec_44_T_3[6:0] ? myVec_53 : _GEN_10846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10848 = 7'h36 == _myNewVec_44_T_3[6:0] ? myVec_54 : _GEN_10847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10849 = 7'h37 == _myNewVec_44_T_3[6:0] ? myVec_55 : _GEN_10848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10850 = 7'h38 == _myNewVec_44_T_3[6:0] ? myVec_56 : _GEN_10849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10851 = 7'h39 == _myNewVec_44_T_3[6:0] ? myVec_57 : _GEN_10850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10852 = 7'h3a == _myNewVec_44_T_3[6:0] ? myVec_58 : _GEN_10851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10853 = 7'h3b == _myNewVec_44_T_3[6:0] ? myVec_59 : _GEN_10852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10854 = 7'h3c == _myNewVec_44_T_3[6:0] ? myVec_60 : _GEN_10853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10855 = 7'h3d == _myNewVec_44_T_3[6:0] ? myVec_61 : _GEN_10854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10856 = 7'h3e == _myNewVec_44_T_3[6:0] ? myVec_62 : _GEN_10855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10857 = 7'h3f == _myNewVec_44_T_3[6:0] ? myVec_63 : _GEN_10856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10858 = 7'h40 == _myNewVec_44_T_3[6:0] ? myVec_64 : _GEN_10857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10859 = 7'h41 == _myNewVec_44_T_3[6:0] ? myVec_65 : _GEN_10858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10860 = 7'h42 == _myNewVec_44_T_3[6:0] ? myVec_66 : _GEN_10859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10861 = 7'h43 == _myNewVec_44_T_3[6:0] ? myVec_67 : _GEN_10860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10862 = 7'h44 == _myNewVec_44_T_3[6:0] ? myVec_68 : _GEN_10861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10863 = 7'h45 == _myNewVec_44_T_3[6:0] ? myVec_69 : _GEN_10862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10864 = 7'h46 == _myNewVec_44_T_3[6:0] ? myVec_70 : _GEN_10863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10865 = 7'h47 == _myNewVec_44_T_3[6:0] ? myVec_71 : _GEN_10864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10866 = 7'h48 == _myNewVec_44_T_3[6:0] ? myVec_72 : _GEN_10865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10867 = 7'h49 == _myNewVec_44_T_3[6:0] ? myVec_73 : _GEN_10866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10868 = 7'h4a == _myNewVec_44_T_3[6:0] ? myVec_74 : _GEN_10867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10869 = 7'h4b == _myNewVec_44_T_3[6:0] ? myVec_75 : _GEN_10868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10870 = 7'h4c == _myNewVec_44_T_3[6:0] ? myVec_76 : _GEN_10869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10871 = 7'h4d == _myNewVec_44_T_3[6:0] ? myVec_77 : _GEN_10870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10872 = 7'h4e == _myNewVec_44_T_3[6:0] ? myVec_78 : _GEN_10871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10873 = 7'h4f == _myNewVec_44_T_3[6:0] ? myVec_79 : _GEN_10872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10874 = 7'h50 == _myNewVec_44_T_3[6:0] ? myVec_80 : _GEN_10873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10875 = 7'h51 == _myNewVec_44_T_3[6:0] ? myVec_81 : _GEN_10874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10876 = 7'h52 == _myNewVec_44_T_3[6:0] ? myVec_82 : _GEN_10875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10877 = 7'h53 == _myNewVec_44_T_3[6:0] ? myVec_83 : _GEN_10876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10878 = 7'h54 == _myNewVec_44_T_3[6:0] ? myVec_84 : _GEN_10877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10879 = 7'h55 == _myNewVec_44_T_3[6:0] ? myVec_85 : _GEN_10878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10880 = 7'h56 == _myNewVec_44_T_3[6:0] ? myVec_86 : _GEN_10879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10881 = 7'h57 == _myNewVec_44_T_3[6:0] ? myVec_87 : _GEN_10880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10882 = 7'h58 == _myNewVec_44_T_3[6:0] ? myVec_88 : _GEN_10881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10883 = 7'h59 == _myNewVec_44_T_3[6:0] ? myVec_89 : _GEN_10882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10884 = 7'h5a == _myNewVec_44_T_3[6:0] ? myVec_90 : _GEN_10883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10885 = 7'h5b == _myNewVec_44_T_3[6:0] ? myVec_91 : _GEN_10884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10886 = 7'h5c == _myNewVec_44_T_3[6:0] ? myVec_92 : _GEN_10885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10887 = 7'h5d == _myNewVec_44_T_3[6:0] ? myVec_93 : _GEN_10886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10888 = 7'h5e == _myNewVec_44_T_3[6:0] ? myVec_94 : _GEN_10887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10889 = 7'h5f == _myNewVec_44_T_3[6:0] ? myVec_95 : _GEN_10888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10890 = 7'h60 == _myNewVec_44_T_3[6:0] ? myVec_96 : _GEN_10889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10891 = 7'h61 == _myNewVec_44_T_3[6:0] ? myVec_97 : _GEN_10890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10892 = 7'h62 == _myNewVec_44_T_3[6:0] ? myVec_98 : _GEN_10891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10893 = 7'h63 == _myNewVec_44_T_3[6:0] ? myVec_99 : _GEN_10892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10894 = 7'h64 == _myNewVec_44_T_3[6:0] ? myVec_100 : _GEN_10893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10895 = 7'h65 == _myNewVec_44_T_3[6:0] ? myVec_101 : _GEN_10894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10896 = 7'h66 == _myNewVec_44_T_3[6:0] ? myVec_102 : _GEN_10895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10897 = 7'h67 == _myNewVec_44_T_3[6:0] ? myVec_103 : _GEN_10896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10898 = 7'h68 == _myNewVec_44_T_3[6:0] ? myVec_104 : _GEN_10897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10899 = 7'h69 == _myNewVec_44_T_3[6:0] ? myVec_105 : _GEN_10898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10900 = 7'h6a == _myNewVec_44_T_3[6:0] ? myVec_106 : _GEN_10899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10901 = 7'h6b == _myNewVec_44_T_3[6:0] ? myVec_107 : _GEN_10900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10902 = 7'h6c == _myNewVec_44_T_3[6:0] ? myVec_108 : _GEN_10901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10903 = 7'h6d == _myNewVec_44_T_3[6:0] ? myVec_109 : _GEN_10902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10904 = 7'h6e == _myNewVec_44_T_3[6:0] ? myVec_110 : _GEN_10903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10905 = 7'h6f == _myNewVec_44_T_3[6:0] ? myVec_111 : _GEN_10904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10906 = 7'h70 == _myNewVec_44_T_3[6:0] ? myVec_112 : _GEN_10905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10907 = 7'h71 == _myNewVec_44_T_3[6:0] ? myVec_113 : _GEN_10906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10908 = 7'h72 == _myNewVec_44_T_3[6:0] ? myVec_114 : _GEN_10907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10909 = 7'h73 == _myNewVec_44_T_3[6:0] ? myVec_115 : _GEN_10908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10910 = 7'h74 == _myNewVec_44_T_3[6:0] ? myVec_116 : _GEN_10909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10911 = 7'h75 == _myNewVec_44_T_3[6:0] ? myVec_117 : _GEN_10910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10912 = 7'h76 == _myNewVec_44_T_3[6:0] ? myVec_118 : _GEN_10911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10913 = 7'h77 == _myNewVec_44_T_3[6:0] ? myVec_119 : _GEN_10912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10914 = 7'h78 == _myNewVec_44_T_3[6:0] ? myVec_120 : _GEN_10913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10915 = 7'h79 == _myNewVec_44_T_3[6:0] ? myVec_121 : _GEN_10914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10916 = 7'h7a == _myNewVec_44_T_3[6:0] ? myVec_122 : _GEN_10915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10917 = 7'h7b == _myNewVec_44_T_3[6:0] ? myVec_123 : _GEN_10916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10918 = 7'h7c == _myNewVec_44_T_3[6:0] ? myVec_124 : _GEN_10917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10919 = 7'h7d == _myNewVec_44_T_3[6:0] ? myVec_125 : _GEN_10918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10920 = 7'h7e == _myNewVec_44_T_3[6:0] ? myVec_126 : _GEN_10919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_44 = 7'h7f == _myNewVec_44_T_3[6:0] ? myVec_127 : _GEN_10920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_43_T_3 = _myNewVec_127_T_1 + 16'h54; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_10923 = 7'h1 == _myNewVec_43_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10924 = 7'h2 == _myNewVec_43_T_3[6:0] ? myVec_2 : _GEN_10923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10925 = 7'h3 == _myNewVec_43_T_3[6:0] ? myVec_3 : _GEN_10924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10926 = 7'h4 == _myNewVec_43_T_3[6:0] ? myVec_4 : _GEN_10925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10927 = 7'h5 == _myNewVec_43_T_3[6:0] ? myVec_5 : _GEN_10926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10928 = 7'h6 == _myNewVec_43_T_3[6:0] ? myVec_6 : _GEN_10927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10929 = 7'h7 == _myNewVec_43_T_3[6:0] ? myVec_7 : _GEN_10928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10930 = 7'h8 == _myNewVec_43_T_3[6:0] ? myVec_8 : _GEN_10929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10931 = 7'h9 == _myNewVec_43_T_3[6:0] ? myVec_9 : _GEN_10930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10932 = 7'ha == _myNewVec_43_T_3[6:0] ? myVec_10 : _GEN_10931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10933 = 7'hb == _myNewVec_43_T_3[6:0] ? myVec_11 : _GEN_10932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10934 = 7'hc == _myNewVec_43_T_3[6:0] ? myVec_12 : _GEN_10933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10935 = 7'hd == _myNewVec_43_T_3[6:0] ? myVec_13 : _GEN_10934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10936 = 7'he == _myNewVec_43_T_3[6:0] ? myVec_14 : _GEN_10935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10937 = 7'hf == _myNewVec_43_T_3[6:0] ? myVec_15 : _GEN_10936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10938 = 7'h10 == _myNewVec_43_T_3[6:0] ? myVec_16 : _GEN_10937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10939 = 7'h11 == _myNewVec_43_T_3[6:0] ? myVec_17 : _GEN_10938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10940 = 7'h12 == _myNewVec_43_T_3[6:0] ? myVec_18 : _GEN_10939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10941 = 7'h13 == _myNewVec_43_T_3[6:0] ? myVec_19 : _GEN_10940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10942 = 7'h14 == _myNewVec_43_T_3[6:0] ? myVec_20 : _GEN_10941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10943 = 7'h15 == _myNewVec_43_T_3[6:0] ? myVec_21 : _GEN_10942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10944 = 7'h16 == _myNewVec_43_T_3[6:0] ? myVec_22 : _GEN_10943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10945 = 7'h17 == _myNewVec_43_T_3[6:0] ? myVec_23 : _GEN_10944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10946 = 7'h18 == _myNewVec_43_T_3[6:0] ? myVec_24 : _GEN_10945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10947 = 7'h19 == _myNewVec_43_T_3[6:0] ? myVec_25 : _GEN_10946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10948 = 7'h1a == _myNewVec_43_T_3[6:0] ? myVec_26 : _GEN_10947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10949 = 7'h1b == _myNewVec_43_T_3[6:0] ? myVec_27 : _GEN_10948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10950 = 7'h1c == _myNewVec_43_T_3[6:0] ? myVec_28 : _GEN_10949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10951 = 7'h1d == _myNewVec_43_T_3[6:0] ? myVec_29 : _GEN_10950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10952 = 7'h1e == _myNewVec_43_T_3[6:0] ? myVec_30 : _GEN_10951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10953 = 7'h1f == _myNewVec_43_T_3[6:0] ? myVec_31 : _GEN_10952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10954 = 7'h20 == _myNewVec_43_T_3[6:0] ? myVec_32 : _GEN_10953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10955 = 7'h21 == _myNewVec_43_T_3[6:0] ? myVec_33 : _GEN_10954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10956 = 7'h22 == _myNewVec_43_T_3[6:0] ? myVec_34 : _GEN_10955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10957 = 7'h23 == _myNewVec_43_T_3[6:0] ? myVec_35 : _GEN_10956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10958 = 7'h24 == _myNewVec_43_T_3[6:0] ? myVec_36 : _GEN_10957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10959 = 7'h25 == _myNewVec_43_T_3[6:0] ? myVec_37 : _GEN_10958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10960 = 7'h26 == _myNewVec_43_T_3[6:0] ? myVec_38 : _GEN_10959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10961 = 7'h27 == _myNewVec_43_T_3[6:0] ? myVec_39 : _GEN_10960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10962 = 7'h28 == _myNewVec_43_T_3[6:0] ? myVec_40 : _GEN_10961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10963 = 7'h29 == _myNewVec_43_T_3[6:0] ? myVec_41 : _GEN_10962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10964 = 7'h2a == _myNewVec_43_T_3[6:0] ? myVec_42 : _GEN_10963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10965 = 7'h2b == _myNewVec_43_T_3[6:0] ? myVec_43 : _GEN_10964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10966 = 7'h2c == _myNewVec_43_T_3[6:0] ? myVec_44 : _GEN_10965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10967 = 7'h2d == _myNewVec_43_T_3[6:0] ? myVec_45 : _GEN_10966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10968 = 7'h2e == _myNewVec_43_T_3[6:0] ? myVec_46 : _GEN_10967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10969 = 7'h2f == _myNewVec_43_T_3[6:0] ? myVec_47 : _GEN_10968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10970 = 7'h30 == _myNewVec_43_T_3[6:0] ? myVec_48 : _GEN_10969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10971 = 7'h31 == _myNewVec_43_T_3[6:0] ? myVec_49 : _GEN_10970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10972 = 7'h32 == _myNewVec_43_T_3[6:0] ? myVec_50 : _GEN_10971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10973 = 7'h33 == _myNewVec_43_T_3[6:0] ? myVec_51 : _GEN_10972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10974 = 7'h34 == _myNewVec_43_T_3[6:0] ? myVec_52 : _GEN_10973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10975 = 7'h35 == _myNewVec_43_T_3[6:0] ? myVec_53 : _GEN_10974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10976 = 7'h36 == _myNewVec_43_T_3[6:0] ? myVec_54 : _GEN_10975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10977 = 7'h37 == _myNewVec_43_T_3[6:0] ? myVec_55 : _GEN_10976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10978 = 7'h38 == _myNewVec_43_T_3[6:0] ? myVec_56 : _GEN_10977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10979 = 7'h39 == _myNewVec_43_T_3[6:0] ? myVec_57 : _GEN_10978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10980 = 7'h3a == _myNewVec_43_T_3[6:0] ? myVec_58 : _GEN_10979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10981 = 7'h3b == _myNewVec_43_T_3[6:0] ? myVec_59 : _GEN_10980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10982 = 7'h3c == _myNewVec_43_T_3[6:0] ? myVec_60 : _GEN_10981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10983 = 7'h3d == _myNewVec_43_T_3[6:0] ? myVec_61 : _GEN_10982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10984 = 7'h3e == _myNewVec_43_T_3[6:0] ? myVec_62 : _GEN_10983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10985 = 7'h3f == _myNewVec_43_T_3[6:0] ? myVec_63 : _GEN_10984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10986 = 7'h40 == _myNewVec_43_T_3[6:0] ? myVec_64 : _GEN_10985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10987 = 7'h41 == _myNewVec_43_T_3[6:0] ? myVec_65 : _GEN_10986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10988 = 7'h42 == _myNewVec_43_T_3[6:0] ? myVec_66 : _GEN_10987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10989 = 7'h43 == _myNewVec_43_T_3[6:0] ? myVec_67 : _GEN_10988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10990 = 7'h44 == _myNewVec_43_T_3[6:0] ? myVec_68 : _GEN_10989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10991 = 7'h45 == _myNewVec_43_T_3[6:0] ? myVec_69 : _GEN_10990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10992 = 7'h46 == _myNewVec_43_T_3[6:0] ? myVec_70 : _GEN_10991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10993 = 7'h47 == _myNewVec_43_T_3[6:0] ? myVec_71 : _GEN_10992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10994 = 7'h48 == _myNewVec_43_T_3[6:0] ? myVec_72 : _GEN_10993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10995 = 7'h49 == _myNewVec_43_T_3[6:0] ? myVec_73 : _GEN_10994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10996 = 7'h4a == _myNewVec_43_T_3[6:0] ? myVec_74 : _GEN_10995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10997 = 7'h4b == _myNewVec_43_T_3[6:0] ? myVec_75 : _GEN_10996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10998 = 7'h4c == _myNewVec_43_T_3[6:0] ? myVec_76 : _GEN_10997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_10999 = 7'h4d == _myNewVec_43_T_3[6:0] ? myVec_77 : _GEN_10998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11000 = 7'h4e == _myNewVec_43_T_3[6:0] ? myVec_78 : _GEN_10999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11001 = 7'h4f == _myNewVec_43_T_3[6:0] ? myVec_79 : _GEN_11000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11002 = 7'h50 == _myNewVec_43_T_3[6:0] ? myVec_80 : _GEN_11001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11003 = 7'h51 == _myNewVec_43_T_3[6:0] ? myVec_81 : _GEN_11002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11004 = 7'h52 == _myNewVec_43_T_3[6:0] ? myVec_82 : _GEN_11003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11005 = 7'h53 == _myNewVec_43_T_3[6:0] ? myVec_83 : _GEN_11004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11006 = 7'h54 == _myNewVec_43_T_3[6:0] ? myVec_84 : _GEN_11005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11007 = 7'h55 == _myNewVec_43_T_3[6:0] ? myVec_85 : _GEN_11006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11008 = 7'h56 == _myNewVec_43_T_3[6:0] ? myVec_86 : _GEN_11007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11009 = 7'h57 == _myNewVec_43_T_3[6:0] ? myVec_87 : _GEN_11008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11010 = 7'h58 == _myNewVec_43_T_3[6:0] ? myVec_88 : _GEN_11009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11011 = 7'h59 == _myNewVec_43_T_3[6:0] ? myVec_89 : _GEN_11010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11012 = 7'h5a == _myNewVec_43_T_3[6:0] ? myVec_90 : _GEN_11011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11013 = 7'h5b == _myNewVec_43_T_3[6:0] ? myVec_91 : _GEN_11012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11014 = 7'h5c == _myNewVec_43_T_3[6:0] ? myVec_92 : _GEN_11013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11015 = 7'h5d == _myNewVec_43_T_3[6:0] ? myVec_93 : _GEN_11014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11016 = 7'h5e == _myNewVec_43_T_3[6:0] ? myVec_94 : _GEN_11015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11017 = 7'h5f == _myNewVec_43_T_3[6:0] ? myVec_95 : _GEN_11016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11018 = 7'h60 == _myNewVec_43_T_3[6:0] ? myVec_96 : _GEN_11017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11019 = 7'h61 == _myNewVec_43_T_3[6:0] ? myVec_97 : _GEN_11018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11020 = 7'h62 == _myNewVec_43_T_3[6:0] ? myVec_98 : _GEN_11019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11021 = 7'h63 == _myNewVec_43_T_3[6:0] ? myVec_99 : _GEN_11020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11022 = 7'h64 == _myNewVec_43_T_3[6:0] ? myVec_100 : _GEN_11021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11023 = 7'h65 == _myNewVec_43_T_3[6:0] ? myVec_101 : _GEN_11022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11024 = 7'h66 == _myNewVec_43_T_3[6:0] ? myVec_102 : _GEN_11023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11025 = 7'h67 == _myNewVec_43_T_3[6:0] ? myVec_103 : _GEN_11024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11026 = 7'h68 == _myNewVec_43_T_3[6:0] ? myVec_104 : _GEN_11025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11027 = 7'h69 == _myNewVec_43_T_3[6:0] ? myVec_105 : _GEN_11026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11028 = 7'h6a == _myNewVec_43_T_3[6:0] ? myVec_106 : _GEN_11027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11029 = 7'h6b == _myNewVec_43_T_3[6:0] ? myVec_107 : _GEN_11028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11030 = 7'h6c == _myNewVec_43_T_3[6:0] ? myVec_108 : _GEN_11029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11031 = 7'h6d == _myNewVec_43_T_3[6:0] ? myVec_109 : _GEN_11030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11032 = 7'h6e == _myNewVec_43_T_3[6:0] ? myVec_110 : _GEN_11031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11033 = 7'h6f == _myNewVec_43_T_3[6:0] ? myVec_111 : _GEN_11032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11034 = 7'h70 == _myNewVec_43_T_3[6:0] ? myVec_112 : _GEN_11033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11035 = 7'h71 == _myNewVec_43_T_3[6:0] ? myVec_113 : _GEN_11034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11036 = 7'h72 == _myNewVec_43_T_3[6:0] ? myVec_114 : _GEN_11035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11037 = 7'h73 == _myNewVec_43_T_3[6:0] ? myVec_115 : _GEN_11036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11038 = 7'h74 == _myNewVec_43_T_3[6:0] ? myVec_116 : _GEN_11037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11039 = 7'h75 == _myNewVec_43_T_3[6:0] ? myVec_117 : _GEN_11038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11040 = 7'h76 == _myNewVec_43_T_3[6:0] ? myVec_118 : _GEN_11039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11041 = 7'h77 == _myNewVec_43_T_3[6:0] ? myVec_119 : _GEN_11040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11042 = 7'h78 == _myNewVec_43_T_3[6:0] ? myVec_120 : _GEN_11041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11043 = 7'h79 == _myNewVec_43_T_3[6:0] ? myVec_121 : _GEN_11042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11044 = 7'h7a == _myNewVec_43_T_3[6:0] ? myVec_122 : _GEN_11043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11045 = 7'h7b == _myNewVec_43_T_3[6:0] ? myVec_123 : _GEN_11044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11046 = 7'h7c == _myNewVec_43_T_3[6:0] ? myVec_124 : _GEN_11045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11047 = 7'h7d == _myNewVec_43_T_3[6:0] ? myVec_125 : _GEN_11046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11048 = 7'h7e == _myNewVec_43_T_3[6:0] ? myVec_126 : _GEN_11047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_43 = 7'h7f == _myNewVec_43_T_3[6:0] ? myVec_127 : _GEN_11048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_42_T_3 = _myNewVec_127_T_1 + 16'h55; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_11051 = 7'h1 == _myNewVec_42_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11052 = 7'h2 == _myNewVec_42_T_3[6:0] ? myVec_2 : _GEN_11051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11053 = 7'h3 == _myNewVec_42_T_3[6:0] ? myVec_3 : _GEN_11052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11054 = 7'h4 == _myNewVec_42_T_3[6:0] ? myVec_4 : _GEN_11053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11055 = 7'h5 == _myNewVec_42_T_3[6:0] ? myVec_5 : _GEN_11054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11056 = 7'h6 == _myNewVec_42_T_3[6:0] ? myVec_6 : _GEN_11055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11057 = 7'h7 == _myNewVec_42_T_3[6:0] ? myVec_7 : _GEN_11056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11058 = 7'h8 == _myNewVec_42_T_3[6:0] ? myVec_8 : _GEN_11057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11059 = 7'h9 == _myNewVec_42_T_3[6:0] ? myVec_9 : _GEN_11058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11060 = 7'ha == _myNewVec_42_T_3[6:0] ? myVec_10 : _GEN_11059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11061 = 7'hb == _myNewVec_42_T_3[6:0] ? myVec_11 : _GEN_11060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11062 = 7'hc == _myNewVec_42_T_3[6:0] ? myVec_12 : _GEN_11061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11063 = 7'hd == _myNewVec_42_T_3[6:0] ? myVec_13 : _GEN_11062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11064 = 7'he == _myNewVec_42_T_3[6:0] ? myVec_14 : _GEN_11063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11065 = 7'hf == _myNewVec_42_T_3[6:0] ? myVec_15 : _GEN_11064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11066 = 7'h10 == _myNewVec_42_T_3[6:0] ? myVec_16 : _GEN_11065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11067 = 7'h11 == _myNewVec_42_T_3[6:0] ? myVec_17 : _GEN_11066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11068 = 7'h12 == _myNewVec_42_T_3[6:0] ? myVec_18 : _GEN_11067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11069 = 7'h13 == _myNewVec_42_T_3[6:0] ? myVec_19 : _GEN_11068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11070 = 7'h14 == _myNewVec_42_T_3[6:0] ? myVec_20 : _GEN_11069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11071 = 7'h15 == _myNewVec_42_T_3[6:0] ? myVec_21 : _GEN_11070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11072 = 7'h16 == _myNewVec_42_T_3[6:0] ? myVec_22 : _GEN_11071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11073 = 7'h17 == _myNewVec_42_T_3[6:0] ? myVec_23 : _GEN_11072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11074 = 7'h18 == _myNewVec_42_T_3[6:0] ? myVec_24 : _GEN_11073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11075 = 7'h19 == _myNewVec_42_T_3[6:0] ? myVec_25 : _GEN_11074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11076 = 7'h1a == _myNewVec_42_T_3[6:0] ? myVec_26 : _GEN_11075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11077 = 7'h1b == _myNewVec_42_T_3[6:0] ? myVec_27 : _GEN_11076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11078 = 7'h1c == _myNewVec_42_T_3[6:0] ? myVec_28 : _GEN_11077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11079 = 7'h1d == _myNewVec_42_T_3[6:0] ? myVec_29 : _GEN_11078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11080 = 7'h1e == _myNewVec_42_T_3[6:0] ? myVec_30 : _GEN_11079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11081 = 7'h1f == _myNewVec_42_T_3[6:0] ? myVec_31 : _GEN_11080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11082 = 7'h20 == _myNewVec_42_T_3[6:0] ? myVec_32 : _GEN_11081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11083 = 7'h21 == _myNewVec_42_T_3[6:0] ? myVec_33 : _GEN_11082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11084 = 7'h22 == _myNewVec_42_T_3[6:0] ? myVec_34 : _GEN_11083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11085 = 7'h23 == _myNewVec_42_T_3[6:0] ? myVec_35 : _GEN_11084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11086 = 7'h24 == _myNewVec_42_T_3[6:0] ? myVec_36 : _GEN_11085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11087 = 7'h25 == _myNewVec_42_T_3[6:0] ? myVec_37 : _GEN_11086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11088 = 7'h26 == _myNewVec_42_T_3[6:0] ? myVec_38 : _GEN_11087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11089 = 7'h27 == _myNewVec_42_T_3[6:0] ? myVec_39 : _GEN_11088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11090 = 7'h28 == _myNewVec_42_T_3[6:0] ? myVec_40 : _GEN_11089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11091 = 7'h29 == _myNewVec_42_T_3[6:0] ? myVec_41 : _GEN_11090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11092 = 7'h2a == _myNewVec_42_T_3[6:0] ? myVec_42 : _GEN_11091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11093 = 7'h2b == _myNewVec_42_T_3[6:0] ? myVec_43 : _GEN_11092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11094 = 7'h2c == _myNewVec_42_T_3[6:0] ? myVec_44 : _GEN_11093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11095 = 7'h2d == _myNewVec_42_T_3[6:0] ? myVec_45 : _GEN_11094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11096 = 7'h2e == _myNewVec_42_T_3[6:0] ? myVec_46 : _GEN_11095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11097 = 7'h2f == _myNewVec_42_T_3[6:0] ? myVec_47 : _GEN_11096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11098 = 7'h30 == _myNewVec_42_T_3[6:0] ? myVec_48 : _GEN_11097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11099 = 7'h31 == _myNewVec_42_T_3[6:0] ? myVec_49 : _GEN_11098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11100 = 7'h32 == _myNewVec_42_T_3[6:0] ? myVec_50 : _GEN_11099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11101 = 7'h33 == _myNewVec_42_T_3[6:0] ? myVec_51 : _GEN_11100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11102 = 7'h34 == _myNewVec_42_T_3[6:0] ? myVec_52 : _GEN_11101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11103 = 7'h35 == _myNewVec_42_T_3[6:0] ? myVec_53 : _GEN_11102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11104 = 7'h36 == _myNewVec_42_T_3[6:0] ? myVec_54 : _GEN_11103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11105 = 7'h37 == _myNewVec_42_T_3[6:0] ? myVec_55 : _GEN_11104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11106 = 7'h38 == _myNewVec_42_T_3[6:0] ? myVec_56 : _GEN_11105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11107 = 7'h39 == _myNewVec_42_T_3[6:0] ? myVec_57 : _GEN_11106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11108 = 7'h3a == _myNewVec_42_T_3[6:0] ? myVec_58 : _GEN_11107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11109 = 7'h3b == _myNewVec_42_T_3[6:0] ? myVec_59 : _GEN_11108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11110 = 7'h3c == _myNewVec_42_T_3[6:0] ? myVec_60 : _GEN_11109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11111 = 7'h3d == _myNewVec_42_T_3[6:0] ? myVec_61 : _GEN_11110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11112 = 7'h3e == _myNewVec_42_T_3[6:0] ? myVec_62 : _GEN_11111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11113 = 7'h3f == _myNewVec_42_T_3[6:0] ? myVec_63 : _GEN_11112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11114 = 7'h40 == _myNewVec_42_T_3[6:0] ? myVec_64 : _GEN_11113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11115 = 7'h41 == _myNewVec_42_T_3[6:0] ? myVec_65 : _GEN_11114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11116 = 7'h42 == _myNewVec_42_T_3[6:0] ? myVec_66 : _GEN_11115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11117 = 7'h43 == _myNewVec_42_T_3[6:0] ? myVec_67 : _GEN_11116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11118 = 7'h44 == _myNewVec_42_T_3[6:0] ? myVec_68 : _GEN_11117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11119 = 7'h45 == _myNewVec_42_T_3[6:0] ? myVec_69 : _GEN_11118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11120 = 7'h46 == _myNewVec_42_T_3[6:0] ? myVec_70 : _GEN_11119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11121 = 7'h47 == _myNewVec_42_T_3[6:0] ? myVec_71 : _GEN_11120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11122 = 7'h48 == _myNewVec_42_T_3[6:0] ? myVec_72 : _GEN_11121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11123 = 7'h49 == _myNewVec_42_T_3[6:0] ? myVec_73 : _GEN_11122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11124 = 7'h4a == _myNewVec_42_T_3[6:0] ? myVec_74 : _GEN_11123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11125 = 7'h4b == _myNewVec_42_T_3[6:0] ? myVec_75 : _GEN_11124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11126 = 7'h4c == _myNewVec_42_T_3[6:0] ? myVec_76 : _GEN_11125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11127 = 7'h4d == _myNewVec_42_T_3[6:0] ? myVec_77 : _GEN_11126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11128 = 7'h4e == _myNewVec_42_T_3[6:0] ? myVec_78 : _GEN_11127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11129 = 7'h4f == _myNewVec_42_T_3[6:0] ? myVec_79 : _GEN_11128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11130 = 7'h50 == _myNewVec_42_T_3[6:0] ? myVec_80 : _GEN_11129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11131 = 7'h51 == _myNewVec_42_T_3[6:0] ? myVec_81 : _GEN_11130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11132 = 7'h52 == _myNewVec_42_T_3[6:0] ? myVec_82 : _GEN_11131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11133 = 7'h53 == _myNewVec_42_T_3[6:0] ? myVec_83 : _GEN_11132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11134 = 7'h54 == _myNewVec_42_T_3[6:0] ? myVec_84 : _GEN_11133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11135 = 7'h55 == _myNewVec_42_T_3[6:0] ? myVec_85 : _GEN_11134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11136 = 7'h56 == _myNewVec_42_T_3[6:0] ? myVec_86 : _GEN_11135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11137 = 7'h57 == _myNewVec_42_T_3[6:0] ? myVec_87 : _GEN_11136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11138 = 7'h58 == _myNewVec_42_T_3[6:0] ? myVec_88 : _GEN_11137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11139 = 7'h59 == _myNewVec_42_T_3[6:0] ? myVec_89 : _GEN_11138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11140 = 7'h5a == _myNewVec_42_T_3[6:0] ? myVec_90 : _GEN_11139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11141 = 7'h5b == _myNewVec_42_T_3[6:0] ? myVec_91 : _GEN_11140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11142 = 7'h5c == _myNewVec_42_T_3[6:0] ? myVec_92 : _GEN_11141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11143 = 7'h5d == _myNewVec_42_T_3[6:0] ? myVec_93 : _GEN_11142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11144 = 7'h5e == _myNewVec_42_T_3[6:0] ? myVec_94 : _GEN_11143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11145 = 7'h5f == _myNewVec_42_T_3[6:0] ? myVec_95 : _GEN_11144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11146 = 7'h60 == _myNewVec_42_T_3[6:0] ? myVec_96 : _GEN_11145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11147 = 7'h61 == _myNewVec_42_T_3[6:0] ? myVec_97 : _GEN_11146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11148 = 7'h62 == _myNewVec_42_T_3[6:0] ? myVec_98 : _GEN_11147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11149 = 7'h63 == _myNewVec_42_T_3[6:0] ? myVec_99 : _GEN_11148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11150 = 7'h64 == _myNewVec_42_T_3[6:0] ? myVec_100 : _GEN_11149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11151 = 7'h65 == _myNewVec_42_T_3[6:0] ? myVec_101 : _GEN_11150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11152 = 7'h66 == _myNewVec_42_T_3[6:0] ? myVec_102 : _GEN_11151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11153 = 7'h67 == _myNewVec_42_T_3[6:0] ? myVec_103 : _GEN_11152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11154 = 7'h68 == _myNewVec_42_T_3[6:0] ? myVec_104 : _GEN_11153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11155 = 7'h69 == _myNewVec_42_T_3[6:0] ? myVec_105 : _GEN_11154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11156 = 7'h6a == _myNewVec_42_T_3[6:0] ? myVec_106 : _GEN_11155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11157 = 7'h6b == _myNewVec_42_T_3[6:0] ? myVec_107 : _GEN_11156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11158 = 7'h6c == _myNewVec_42_T_3[6:0] ? myVec_108 : _GEN_11157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11159 = 7'h6d == _myNewVec_42_T_3[6:0] ? myVec_109 : _GEN_11158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11160 = 7'h6e == _myNewVec_42_T_3[6:0] ? myVec_110 : _GEN_11159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11161 = 7'h6f == _myNewVec_42_T_3[6:0] ? myVec_111 : _GEN_11160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11162 = 7'h70 == _myNewVec_42_T_3[6:0] ? myVec_112 : _GEN_11161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11163 = 7'h71 == _myNewVec_42_T_3[6:0] ? myVec_113 : _GEN_11162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11164 = 7'h72 == _myNewVec_42_T_3[6:0] ? myVec_114 : _GEN_11163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11165 = 7'h73 == _myNewVec_42_T_3[6:0] ? myVec_115 : _GEN_11164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11166 = 7'h74 == _myNewVec_42_T_3[6:0] ? myVec_116 : _GEN_11165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11167 = 7'h75 == _myNewVec_42_T_3[6:0] ? myVec_117 : _GEN_11166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11168 = 7'h76 == _myNewVec_42_T_3[6:0] ? myVec_118 : _GEN_11167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11169 = 7'h77 == _myNewVec_42_T_3[6:0] ? myVec_119 : _GEN_11168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11170 = 7'h78 == _myNewVec_42_T_3[6:0] ? myVec_120 : _GEN_11169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11171 = 7'h79 == _myNewVec_42_T_3[6:0] ? myVec_121 : _GEN_11170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11172 = 7'h7a == _myNewVec_42_T_3[6:0] ? myVec_122 : _GEN_11171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11173 = 7'h7b == _myNewVec_42_T_3[6:0] ? myVec_123 : _GEN_11172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11174 = 7'h7c == _myNewVec_42_T_3[6:0] ? myVec_124 : _GEN_11173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11175 = 7'h7d == _myNewVec_42_T_3[6:0] ? myVec_125 : _GEN_11174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11176 = 7'h7e == _myNewVec_42_T_3[6:0] ? myVec_126 : _GEN_11175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_42 = 7'h7f == _myNewVec_42_T_3[6:0] ? myVec_127 : _GEN_11176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_41_T_3 = _myNewVec_127_T_1 + 16'h56; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_11179 = 7'h1 == _myNewVec_41_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11180 = 7'h2 == _myNewVec_41_T_3[6:0] ? myVec_2 : _GEN_11179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11181 = 7'h3 == _myNewVec_41_T_3[6:0] ? myVec_3 : _GEN_11180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11182 = 7'h4 == _myNewVec_41_T_3[6:0] ? myVec_4 : _GEN_11181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11183 = 7'h5 == _myNewVec_41_T_3[6:0] ? myVec_5 : _GEN_11182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11184 = 7'h6 == _myNewVec_41_T_3[6:0] ? myVec_6 : _GEN_11183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11185 = 7'h7 == _myNewVec_41_T_3[6:0] ? myVec_7 : _GEN_11184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11186 = 7'h8 == _myNewVec_41_T_3[6:0] ? myVec_8 : _GEN_11185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11187 = 7'h9 == _myNewVec_41_T_3[6:0] ? myVec_9 : _GEN_11186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11188 = 7'ha == _myNewVec_41_T_3[6:0] ? myVec_10 : _GEN_11187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11189 = 7'hb == _myNewVec_41_T_3[6:0] ? myVec_11 : _GEN_11188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11190 = 7'hc == _myNewVec_41_T_3[6:0] ? myVec_12 : _GEN_11189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11191 = 7'hd == _myNewVec_41_T_3[6:0] ? myVec_13 : _GEN_11190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11192 = 7'he == _myNewVec_41_T_3[6:0] ? myVec_14 : _GEN_11191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11193 = 7'hf == _myNewVec_41_T_3[6:0] ? myVec_15 : _GEN_11192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11194 = 7'h10 == _myNewVec_41_T_3[6:0] ? myVec_16 : _GEN_11193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11195 = 7'h11 == _myNewVec_41_T_3[6:0] ? myVec_17 : _GEN_11194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11196 = 7'h12 == _myNewVec_41_T_3[6:0] ? myVec_18 : _GEN_11195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11197 = 7'h13 == _myNewVec_41_T_3[6:0] ? myVec_19 : _GEN_11196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11198 = 7'h14 == _myNewVec_41_T_3[6:0] ? myVec_20 : _GEN_11197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11199 = 7'h15 == _myNewVec_41_T_3[6:0] ? myVec_21 : _GEN_11198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11200 = 7'h16 == _myNewVec_41_T_3[6:0] ? myVec_22 : _GEN_11199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11201 = 7'h17 == _myNewVec_41_T_3[6:0] ? myVec_23 : _GEN_11200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11202 = 7'h18 == _myNewVec_41_T_3[6:0] ? myVec_24 : _GEN_11201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11203 = 7'h19 == _myNewVec_41_T_3[6:0] ? myVec_25 : _GEN_11202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11204 = 7'h1a == _myNewVec_41_T_3[6:0] ? myVec_26 : _GEN_11203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11205 = 7'h1b == _myNewVec_41_T_3[6:0] ? myVec_27 : _GEN_11204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11206 = 7'h1c == _myNewVec_41_T_3[6:0] ? myVec_28 : _GEN_11205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11207 = 7'h1d == _myNewVec_41_T_3[6:0] ? myVec_29 : _GEN_11206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11208 = 7'h1e == _myNewVec_41_T_3[6:0] ? myVec_30 : _GEN_11207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11209 = 7'h1f == _myNewVec_41_T_3[6:0] ? myVec_31 : _GEN_11208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11210 = 7'h20 == _myNewVec_41_T_3[6:0] ? myVec_32 : _GEN_11209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11211 = 7'h21 == _myNewVec_41_T_3[6:0] ? myVec_33 : _GEN_11210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11212 = 7'h22 == _myNewVec_41_T_3[6:0] ? myVec_34 : _GEN_11211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11213 = 7'h23 == _myNewVec_41_T_3[6:0] ? myVec_35 : _GEN_11212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11214 = 7'h24 == _myNewVec_41_T_3[6:0] ? myVec_36 : _GEN_11213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11215 = 7'h25 == _myNewVec_41_T_3[6:0] ? myVec_37 : _GEN_11214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11216 = 7'h26 == _myNewVec_41_T_3[6:0] ? myVec_38 : _GEN_11215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11217 = 7'h27 == _myNewVec_41_T_3[6:0] ? myVec_39 : _GEN_11216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11218 = 7'h28 == _myNewVec_41_T_3[6:0] ? myVec_40 : _GEN_11217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11219 = 7'h29 == _myNewVec_41_T_3[6:0] ? myVec_41 : _GEN_11218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11220 = 7'h2a == _myNewVec_41_T_3[6:0] ? myVec_42 : _GEN_11219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11221 = 7'h2b == _myNewVec_41_T_3[6:0] ? myVec_43 : _GEN_11220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11222 = 7'h2c == _myNewVec_41_T_3[6:0] ? myVec_44 : _GEN_11221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11223 = 7'h2d == _myNewVec_41_T_3[6:0] ? myVec_45 : _GEN_11222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11224 = 7'h2e == _myNewVec_41_T_3[6:0] ? myVec_46 : _GEN_11223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11225 = 7'h2f == _myNewVec_41_T_3[6:0] ? myVec_47 : _GEN_11224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11226 = 7'h30 == _myNewVec_41_T_3[6:0] ? myVec_48 : _GEN_11225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11227 = 7'h31 == _myNewVec_41_T_3[6:0] ? myVec_49 : _GEN_11226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11228 = 7'h32 == _myNewVec_41_T_3[6:0] ? myVec_50 : _GEN_11227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11229 = 7'h33 == _myNewVec_41_T_3[6:0] ? myVec_51 : _GEN_11228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11230 = 7'h34 == _myNewVec_41_T_3[6:0] ? myVec_52 : _GEN_11229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11231 = 7'h35 == _myNewVec_41_T_3[6:0] ? myVec_53 : _GEN_11230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11232 = 7'h36 == _myNewVec_41_T_3[6:0] ? myVec_54 : _GEN_11231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11233 = 7'h37 == _myNewVec_41_T_3[6:0] ? myVec_55 : _GEN_11232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11234 = 7'h38 == _myNewVec_41_T_3[6:0] ? myVec_56 : _GEN_11233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11235 = 7'h39 == _myNewVec_41_T_3[6:0] ? myVec_57 : _GEN_11234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11236 = 7'h3a == _myNewVec_41_T_3[6:0] ? myVec_58 : _GEN_11235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11237 = 7'h3b == _myNewVec_41_T_3[6:0] ? myVec_59 : _GEN_11236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11238 = 7'h3c == _myNewVec_41_T_3[6:0] ? myVec_60 : _GEN_11237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11239 = 7'h3d == _myNewVec_41_T_3[6:0] ? myVec_61 : _GEN_11238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11240 = 7'h3e == _myNewVec_41_T_3[6:0] ? myVec_62 : _GEN_11239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11241 = 7'h3f == _myNewVec_41_T_3[6:0] ? myVec_63 : _GEN_11240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11242 = 7'h40 == _myNewVec_41_T_3[6:0] ? myVec_64 : _GEN_11241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11243 = 7'h41 == _myNewVec_41_T_3[6:0] ? myVec_65 : _GEN_11242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11244 = 7'h42 == _myNewVec_41_T_3[6:0] ? myVec_66 : _GEN_11243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11245 = 7'h43 == _myNewVec_41_T_3[6:0] ? myVec_67 : _GEN_11244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11246 = 7'h44 == _myNewVec_41_T_3[6:0] ? myVec_68 : _GEN_11245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11247 = 7'h45 == _myNewVec_41_T_3[6:0] ? myVec_69 : _GEN_11246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11248 = 7'h46 == _myNewVec_41_T_3[6:0] ? myVec_70 : _GEN_11247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11249 = 7'h47 == _myNewVec_41_T_3[6:0] ? myVec_71 : _GEN_11248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11250 = 7'h48 == _myNewVec_41_T_3[6:0] ? myVec_72 : _GEN_11249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11251 = 7'h49 == _myNewVec_41_T_3[6:0] ? myVec_73 : _GEN_11250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11252 = 7'h4a == _myNewVec_41_T_3[6:0] ? myVec_74 : _GEN_11251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11253 = 7'h4b == _myNewVec_41_T_3[6:0] ? myVec_75 : _GEN_11252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11254 = 7'h4c == _myNewVec_41_T_3[6:0] ? myVec_76 : _GEN_11253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11255 = 7'h4d == _myNewVec_41_T_3[6:0] ? myVec_77 : _GEN_11254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11256 = 7'h4e == _myNewVec_41_T_3[6:0] ? myVec_78 : _GEN_11255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11257 = 7'h4f == _myNewVec_41_T_3[6:0] ? myVec_79 : _GEN_11256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11258 = 7'h50 == _myNewVec_41_T_3[6:0] ? myVec_80 : _GEN_11257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11259 = 7'h51 == _myNewVec_41_T_3[6:0] ? myVec_81 : _GEN_11258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11260 = 7'h52 == _myNewVec_41_T_3[6:0] ? myVec_82 : _GEN_11259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11261 = 7'h53 == _myNewVec_41_T_3[6:0] ? myVec_83 : _GEN_11260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11262 = 7'h54 == _myNewVec_41_T_3[6:0] ? myVec_84 : _GEN_11261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11263 = 7'h55 == _myNewVec_41_T_3[6:0] ? myVec_85 : _GEN_11262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11264 = 7'h56 == _myNewVec_41_T_3[6:0] ? myVec_86 : _GEN_11263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11265 = 7'h57 == _myNewVec_41_T_3[6:0] ? myVec_87 : _GEN_11264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11266 = 7'h58 == _myNewVec_41_T_3[6:0] ? myVec_88 : _GEN_11265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11267 = 7'h59 == _myNewVec_41_T_3[6:0] ? myVec_89 : _GEN_11266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11268 = 7'h5a == _myNewVec_41_T_3[6:0] ? myVec_90 : _GEN_11267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11269 = 7'h5b == _myNewVec_41_T_3[6:0] ? myVec_91 : _GEN_11268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11270 = 7'h5c == _myNewVec_41_T_3[6:0] ? myVec_92 : _GEN_11269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11271 = 7'h5d == _myNewVec_41_T_3[6:0] ? myVec_93 : _GEN_11270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11272 = 7'h5e == _myNewVec_41_T_3[6:0] ? myVec_94 : _GEN_11271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11273 = 7'h5f == _myNewVec_41_T_3[6:0] ? myVec_95 : _GEN_11272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11274 = 7'h60 == _myNewVec_41_T_3[6:0] ? myVec_96 : _GEN_11273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11275 = 7'h61 == _myNewVec_41_T_3[6:0] ? myVec_97 : _GEN_11274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11276 = 7'h62 == _myNewVec_41_T_3[6:0] ? myVec_98 : _GEN_11275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11277 = 7'h63 == _myNewVec_41_T_3[6:0] ? myVec_99 : _GEN_11276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11278 = 7'h64 == _myNewVec_41_T_3[6:0] ? myVec_100 : _GEN_11277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11279 = 7'h65 == _myNewVec_41_T_3[6:0] ? myVec_101 : _GEN_11278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11280 = 7'h66 == _myNewVec_41_T_3[6:0] ? myVec_102 : _GEN_11279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11281 = 7'h67 == _myNewVec_41_T_3[6:0] ? myVec_103 : _GEN_11280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11282 = 7'h68 == _myNewVec_41_T_3[6:0] ? myVec_104 : _GEN_11281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11283 = 7'h69 == _myNewVec_41_T_3[6:0] ? myVec_105 : _GEN_11282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11284 = 7'h6a == _myNewVec_41_T_3[6:0] ? myVec_106 : _GEN_11283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11285 = 7'h6b == _myNewVec_41_T_3[6:0] ? myVec_107 : _GEN_11284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11286 = 7'h6c == _myNewVec_41_T_3[6:0] ? myVec_108 : _GEN_11285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11287 = 7'h6d == _myNewVec_41_T_3[6:0] ? myVec_109 : _GEN_11286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11288 = 7'h6e == _myNewVec_41_T_3[6:0] ? myVec_110 : _GEN_11287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11289 = 7'h6f == _myNewVec_41_T_3[6:0] ? myVec_111 : _GEN_11288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11290 = 7'h70 == _myNewVec_41_T_3[6:0] ? myVec_112 : _GEN_11289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11291 = 7'h71 == _myNewVec_41_T_3[6:0] ? myVec_113 : _GEN_11290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11292 = 7'h72 == _myNewVec_41_T_3[6:0] ? myVec_114 : _GEN_11291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11293 = 7'h73 == _myNewVec_41_T_3[6:0] ? myVec_115 : _GEN_11292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11294 = 7'h74 == _myNewVec_41_T_3[6:0] ? myVec_116 : _GEN_11293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11295 = 7'h75 == _myNewVec_41_T_3[6:0] ? myVec_117 : _GEN_11294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11296 = 7'h76 == _myNewVec_41_T_3[6:0] ? myVec_118 : _GEN_11295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11297 = 7'h77 == _myNewVec_41_T_3[6:0] ? myVec_119 : _GEN_11296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11298 = 7'h78 == _myNewVec_41_T_3[6:0] ? myVec_120 : _GEN_11297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11299 = 7'h79 == _myNewVec_41_T_3[6:0] ? myVec_121 : _GEN_11298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11300 = 7'h7a == _myNewVec_41_T_3[6:0] ? myVec_122 : _GEN_11299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11301 = 7'h7b == _myNewVec_41_T_3[6:0] ? myVec_123 : _GEN_11300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11302 = 7'h7c == _myNewVec_41_T_3[6:0] ? myVec_124 : _GEN_11301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11303 = 7'h7d == _myNewVec_41_T_3[6:0] ? myVec_125 : _GEN_11302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11304 = 7'h7e == _myNewVec_41_T_3[6:0] ? myVec_126 : _GEN_11303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_41 = 7'h7f == _myNewVec_41_T_3[6:0] ? myVec_127 : _GEN_11304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_40_T_3 = _myNewVec_127_T_1 + 16'h57; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_11307 = 7'h1 == _myNewVec_40_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11308 = 7'h2 == _myNewVec_40_T_3[6:0] ? myVec_2 : _GEN_11307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11309 = 7'h3 == _myNewVec_40_T_3[6:0] ? myVec_3 : _GEN_11308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11310 = 7'h4 == _myNewVec_40_T_3[6:0] ? myVec_4 : _GEN_11309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11311 = 7'h5 == _myNewVec_40_T_3[6:0] ? myVec_5 : _GEN_11310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11312 = 7'h6 == _myNewVec_40_T_3[6:0] ? myVec_6 : _GEN_11311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11313 = 7'h7 == _myNewVec_40_T_3[6:0] ? myVec_7 : _GEN_11312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11314 = 7'h8 == _myNewVec_40_T_3[6:0] ? myVec_8 : _GEN_11313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11315 = 7'h9 == _myNewVec_40_T_3[6:0] ? myVec_9 : _GEN_11314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11316 = 7'ha == _myNewVec_40_T_3[6:0] ? myVec_10 : _GEN_11315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11317 = 7'hb == _myNewVec_40_T_3[6:0] ? myVec_11 : _GEN_11316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11318 = 7'hc == _myNewVec_40_T_3[6:0] ? myVec_12 : _GEN_11317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11319 = 7'hd == _myNewVec_40_T_3[6:0] ? myVec_13 : _GEN_11318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11320 = 7'he == _myNewVec_40_T_3[6:0] ? myVec_14 : _GEN_11319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11321 = 7'hf == _myNewVec_40_T_3[6:0] ? myVec_15 : _GEN_11320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11322 = 7'h10 == _myNewVec_40_T_3[6:0] ? myVec_16 : _GEN_11321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11323 = 7'h11 == _myNewVec_40_T_3[6:0] ? myVec_17 : _GEN_11322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11324 = 7'h12 == _myNewVec_40_T_3[6:0] ? myVec_18 : _GEN_11323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11325 = 7'h13 == _myNewVec_40_T_3[6:0] ? myVec_19 : _GEN_11324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11326 = 7'h14 == _myNewVec_40_T_3[6:0] ? myVec_20 : _GEN_11325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11327 = 7'h15 == _myNewVec_40_T_3[6:0] ? myVec_21 : _GEN_11326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11328 = 7'h16 == _myNewVec_40_T_3[6:0] ? myVec_22 : _GEN_11327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11329 = 7'h17 == _myNewVec_40_T_3[6:0] ? myVec_23 : _GEN_11328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11330 = 7'h18 == _myNewVec_40_T_3[6:0] ? myVec_24 : _GEN_11329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11331 = 7'h19 == _myNewVec_40_T_3[6:0] ? myVec_25 : _GEN_11330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11332 = 7'h1a == _myNewVec_40_T_3[6:0] ? myVec_26 : _GEN_11331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11333 = 7'h1b == _myNewVec_40_T_3[6:0] ? myVec_27 : _GEN_11332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11334 = 7'h1c == _myNewVec_40_T_3[6:0] ? myVec_28 : _GEN_11333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11335 = 7'h1d == _myNewVec_40_T_3[6:0] ? myVec_29 : _GEN_11334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11336 = 7'h1e == _myNewVec_40_T_3[6:0] ? myVec_30 : _GEN_11335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11337 = 7'h1f == _myNewVec_40_T_3[6:0] ? myVec_31 : _GEN_11336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11338 = 7'h20 == _myNewVec_40_T_3[6:0] ? myVec_32 : _GEN_11337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11339 = 7'h21 == _myNewVec_40_T_3[6:0] ? myVec_33 : _GEN_11338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11340 = 7'h22 == _myNewVec_40_T_3[6:0] ? myVec_34 : _GEN_11339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11341 = 7'h23 == _myNewVec_40_T_3[6:0] ? myVec_35 : _GEN_11340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11342 = 7'h24 == _myNewVec_40_T_3[6:0] ? myVec_36 : _GEN_11341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11343 = 7'h25 == _myNewVec_40_T_3[6:0] ? myVec_37 : _GEN_11342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11344 = 7'h26 == _myNewVec_40_T_3[6:0] ? myVec_38 : _GEN_11343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11345 = 7'h27 == _myNewVec_40_T_3[6:0] ? myVec_39 : _GEN_11344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11346 = 7'h28 == _myNewVec_40_T_3[6:0] ? myVec_40 : _GEN_11345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11347 = 7'h29 == _myNewVec_40_T_3[6:0] ? myVec_41 : _GEN_11346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11348 = 7'h2a == _myNewVec_40_T_3[6:0] ? myVec_42 : _GEN_11347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11349 = 7'h2b == _myNewVec_40_T_3[6:0] ? myVec_43 : _GEN_11348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11350 = 7'h2c == _myNewVec_40_T_3[6:0] ? myVec_44 : _GEN_11349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11351 = 7'h2d == _myNewVec_40_T_3[6:0] ? myVec_45 : _GEN_11350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11352 = 7'h2e == _myNewVec_40_T_3[6:0] ? myVec_46 : _GEN_11351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11353 = 7'h2f == _myNewVec_40_T_3[6:0] ? myVec_47 : _GEN_11352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11354 = 7'h30 == _myNewVec_40_T_3[6:0] ? myVec_48 : _GEN_11353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11355 = 7'h31 == _myNewVec_40_T_3[6:0] ? myVec_49 : _GEN_11354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11356 = 7'h32 == _myNewVec_40_T_3[6:0] ? myVec_50 : _GEN_11355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11357 = 7'h33 == _myNewVec_40_T_3[6:0] ? myVec_51 : _GEN_11356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11358 = 7'h34 == _myNewVec_40_T_3[6:0] ? myVec_52 : _GEN_11357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11359 = 7'h35 == _myNewVec_40_T_3[6:0] ? myVec_53 : _GEN_11358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11360 = 7'h36 == _myNewVec_40_T_3[6:0] ? myVec_54 : _GEN_11359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11361 = 7'h37 == _myNewVec_40_T_3[6:0] ? myVec_55 : _GEN_11360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11362 = 7'h38 == _myNewVec_40_T_3[6:0] ? myVec_56 : _GEN_11361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11363 = 7'h39 == _myNewVec_40_T_3[6:0] ? myVec_57 : _GEN_11362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11364 = 7'h3a == _myNewVec_40_T_3[6:0] ? myVec_58 : _GEN_11363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11365 = 7'h3b == _myNewVec_40_T_3[6:0] ? myVec_59 : _GEN_11364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11366 = 7'h3c == _myNewVec_40_T_3[6:0] ? myVec_60 : _GEN_11365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11367 = 7'h3d == _myNewVec_40_T_3[6:0] ? myVec_61 : _GEN_11366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11368 = 7'h3e == _myNewVec_40_T_3[6:0] ? myVec_62 : _GEN_11367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11369 = 7'h3f == _myNewVec_40_T_3[6:0] ? myVec_63 : _GEN_11368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11370 = 7'h40 == _myNewVec_40_T_3[6:0] ? myVec_64 : _GEN_11369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11371 = 7'h41 == _myNewVec_40_T_3[6:0] ? myVec_65 : _GEN_11370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11372 = 7'h42 == _myNewVec_40_T_3[6:0] ? myVec_66 : _GEN_11371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11373 = 7'h43 == _myNewVec_40_T_3[6:0] ? myVec_67 : _GEN_11372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11374 = 7'h44 == _myNewVec_40_T_3[6:0] ? myVec_68 : _GEN_11373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11375 = 7'h45 == _myNewVec_40_T_3[6:0] ? myVec_69 : _GEN_11374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11376 = 7'h46 == _myNewVec_40_T_3[6:0] ? myVec_70 : _GEN_11375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11377 = 7'h47 == _myNewVec_40_T_3[6:0] ? myVec_71 : _GEN_11376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11378 = 7'h48 == _myNewVec_40_T_3[6:0] ? myVec_72 : _GEN_11377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11379 = 7'h49 == _myNewVec_40_T_3[6:0] ? myVec_73 : _GEN_11378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11380 = 7'h4a == _myNewVec_40_T_3[6:0] ? myVec_74 : _GEN_11379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11381 = 7'h4b == _myNewVec_40_T_3[6:0] ? myVec_75 : _GEN_11380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11382 = 7'h4c == _myNewVec_40_T_3[6:0] ? myVec_76 : _GEN_11381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11383 = 7'h4d == _myNewVec_40_T_3[6:0] ? myVec_77 : _GEN_11382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11384 = 7'h4e == _myNewVec_40_T_3[6:0] ? myVec_78 : _GEN_11383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11385 = 7'h4f == _myNewVec_40_T_3[6:0] ? myVec_79 : _GEN_11384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11386 = 7'h50 == _myNewVec_40_T_3[6:0] ? myVec_80 : _GEN_11385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11387 = 7'h51 == _myNewVec_40_T_3[6:0] ? myVec_81 : _GEN_11386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11388 = 7'h52 == _myNewVec_40_T_3[6:0] ? myVec_82 : _GEN_11387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11389 = 7'h53 == _myNewVec_40_T_3[6:0] ? myVec_83 : _GEN_11388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11390 = 7'h54 == _myNewVec_40_T_3[6:0] ? myVec_84 : _GEN_11389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11391 = 7'h55 == _myNewVec_40_T_3[6:0] ? myVec_85 : _GEN_11390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11392 = 7'h56 == _myNewVec_40_T_3[6:0] ? myVec_86 : _GEN_11391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11393 = 7'h57 == _myNewVec_40_T_3[6:0] ? myVec_87 : _GEN_11392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11394 = 7'h58 == _myNewVec_40_T_3[6:0] ? myVec_88 : _GEN_11393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11395 = 7'h59 == _myNewVec_40_T_3[6:0] ? myVec_89 : _GEN_11394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11396 = 7'h5a == _myNewVec_40_T_3[6:0] ? myVec_90 : _GEN_11395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11397 = 7'h5b == _myNewVec_40_T_3[6:0] ? myVec_91 : _GEN_11396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11398 = 7'h5c == _myNewVec_40_T_3[6:0] ? myVec_92 : _GEN_11397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11399 = 7'h5d == _myNewVec_40_T_3[6:0] ? myVec_93 : _GEN_11398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11400 = 7'h5e == _myNewVec_40_T_3[6:0] ? myVec_94 : _GEN_11399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11401 = 7'h5f == _myNewVec_40_T_3[6:0] ? myVec_95 : _GEN_11400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11402 = 7'h60 == _myNewVec_40_T_3[6:0] ? myVec_96 : _GEN_11401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11403 = 7'h61 == _myNewVec_40_T_3[6:0] ? myVec_97 : _GEN_11402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11404 = 7'h62 == _myNewVec_40_T_3[6:0] ? myVec_98 : _GEN_11403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11405 = 7'h63 == _myNewVec_40_T_3[6:0] ? myVec_99 : _GEN_11404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11406 = 7'h64 == _myNewVec_40_T_3[6:0] ? myVec_100 : _GEN_11405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11407 = 7'h65 == _myNewVec_40_T_3[6:0] ? myVec_101 : _GEN_11406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11408 = 7'h66 == _myNewVec_40_T_3[6:0] ? myVec_102 : _GEN_11407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11409 = 7'h67 == _myNewVec_40_T_3[6:0] ? myVec_103 : _GEN_11408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11410 = 7'h68 == _myNewVec_40_T_3[6:0] ? myVec_104 : _GEN_11409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11411 = 7'h69 == _myNewVec_40_T_3[6:0] ? myVec_105 : _GEN_11410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11412 = 7'h6a == _myNewVec_40_T_3[6:0] ? myVec_106 : _GEN_11411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11413 = 7'h6b == _myNewVec_40_T_3[6:0] ? myVec_107 : _GEN_11412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11414 = 7'h6c == _myNewVec_40_T_3[6:0] ? myVec_108 : _GEN_11413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11415 = 7'h6d == _myNewVec_40_T_3[6:0] ? myVec_109 : _GEN_11414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11416 = 7'h6e == _myNewVec_40_T_3[6:0] ? myVec_110 : _GEN_11415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11417 = 7'h6f == _myNewVec_40_T_3[6:0] ? myVec_111 : _GEN_11416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11418 = 7'h70 == _myNewVec_40_T_3[6:0] ? myVec_112 : _GEN_11417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11419 = 7'h71 == _myNewVec_40_T_3[6:0] ? myVec_113 : _GEN_11418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11420 = 7'h72 == _myNewVec_40_T_3[6:0] ? myVec_114 : _GEN_11419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11421 = 7'h73 == _myNewVec_40_T_3[6:0] ? myVec_115 : _GEN_11420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11422 = 7'h74 == _myNewVec_40_T_3[6:0] ? myVec_116 : _GEN_11421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11423 = 7'h75 == _myNewVec_40_T_3[6:0] ? myVec_117 : _GEN_11422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11424 = 7'h76 == _myNewVec_40_T_3[6:0] ? myVec_118 : _GEN_11423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11425 = 7'h77 == _myNewVec_40_T_3[6:0] ? myVec_119 : _GEN_11424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11426 = 7'h78 == _myNewVec_40_T_3[6:0] ? myVec_120 : _GEN_11425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11427 = 7'h79 == _myNewVec_40_T_3[6:0] ? myVec_121 : _GEN_11426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11428 = 7'h7a == _myNewVec_40_T_3[6:0] ? myVec_122 : _GEN_11427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11429 = 7'h7b == _myNewVec_40_T_3[6:0] ? myVec_123 : _GEN_11428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11430 = 7'h7c == _myNewVec_40_T_3[6:0] ? myVec_124 : _GEN_11429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11431 = 7'h7d == _myNewVec_40_T_3[6:0] ? myVec_125 : _GEN_11430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11432 = 7'h7e == _myNewVec_40_T_3[6:0] ? myVec_126 : _GEN_11431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_40 = 7'h7f == _myNewVec_40_T_3[6:0] ? myVec_127 : _GEN_11432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_39_T_3 = _myNewVec_127_T_1 + 16'h58; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_11435 = 7'h1 == _myNewVec_39_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11436 = 7'h2 == _myNewVec_39_T_3[6:0] ? myVec_2 : _GEN_11435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11437 = 7'h3 == _myNewVec_39_T_3[6:0] ? myVec_3 : _GEN_11436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11438 = 7'h4 == _myNewVec_39_T_3[6:0] ? myVec_4 : _GEN_11437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11439 = 7'h5 == _myNewVec_39_T_3[6:0] ? myVec_5 : _GEN_11438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11440 = 7'h6 == _myNewVec_39_T_3[6:0] ? myVec_6 : _GEN_11439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11441 = 7'h7 == _myNewVec_39_T_3[6:0] ? myVec_7 : _GEN_11440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11442 = 7'h8 == _myNewVec_39_T_3[6:0] ? myVec_8 : _GEN_11441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11443 = 7'h9 == _myNewVec_39_T_3[6:0] ? myVec_9 : _GEN_11442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11444 = 7'ha == _myNewVec_39_T_3[6:0] ? myVec_10 : _GEN_11443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11445 = 7'hb == _myNewVec_39_T_3[6:0] ? myVec_11 : _GEN_11444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11446 = 7'hc == _myNewVec_39_T_3[6:0] ? myVec_12 : _GEN_11445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11447 = 7'hd == _myNewVec_39_T_3[6:0] ? myVec_13 : _GEN_11446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11448 = 7'he == _myNewVec_39_T_3[6:0] ? myVec_14 : _GEN_11447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11449 = 7'hf == _myNewVec_39_T_3[6:0] ? myVec_15 : _GEN_11448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11450 = 7'h10 == _myNewVec_39_T_3[6:0] ? myVec_16 : _GEN_11449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11451 = 7'h11 == _myNewVec_39_T_3[6:0] ? myVec_17 : _GEN_11450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11452 = 7'h12 == _myNewVec_39_T_3[6:0] ? myVec_18 : _GEN_11451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11453 = 7'h13 == _myNewVec_39_T_3[6:0] ? myVec_19 : _GEN_11452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11454 = 7'h14 == _myNewVec_39_T_3[6:0] ? myVec_20 : _GEN_11453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11455 = 7'h15 == _myNewVec_39_T_3[6:0] ? myVec_21 : _GEN_11454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11456 = 7'h16 == _myNewVec_39_T_3[6:0] ? myVec_22 : _GEN_11455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11457 = 7'h17 == _myNewVec_39_T_3[6:0] ? myVec_23 : _GEN_11456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11458 = 7'h18 == _myNewVec_39_T_3[6:0] ? myVec_24 : _GEN_11457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11459 = 7'h19 == _myNewVec_39_T_3[6:0] ? myVec_25 : _GEN_11458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11460 = 7'h1a == _myNewVec_39_T_3[6:0] ? myVec_26 : _GEN_11459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11461 = 7'h1b == _myNewVec_39_T_3[6:0] ? myVec_27 : _GEN_11460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11462 = 7'h1c == _myNewVec_39_T_3[6:0] ? myVec_28 : _GEN_11461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11463 = 7'h1d == _myNewVec_39_T_3[6:0] ? myVec_29 : _GEN_11462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11464 = 7'h1e == _myNewVec_39_T_3[6:0] ? myVec_30 : _GEN_11463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11465 = 7'h1f == _myNewVec_39_T_3[6:0] ? myVec_31 : _GEN_11464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11466 = 7'h20 == _myNewVec_39_T_3[6:0] ? myVec_32 : _GEN_11465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11467 = 7'h21 == _myNewVec_39_T_3[6:0] ? myVec_33 : _GEN_11466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11468 = 7'h22 == _myNewVec_39_T_3[6:0] ? myVec_34 : _GEN_11467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11469 = 7'h23 == _myNewVec_39_T_3[6:0] ? myVec_35 : _GEN_11468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11470 = 7'h24 == _myNewVec_39_T_3[6:0] ? myVec_36 : _GEN_11469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11471 = 7'h25 == _myNewVec_39_T_3[6:0] ? myVec_37 : _GEN_11470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11472 = 7'h26 == _myNewVec_39_T_3[6:0] ? myVec_38 : _GEN_11471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11473 = 7'h27 == _myNewVec_39_T_3[6:0] ? myVec_39 : _GEN_11472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11474 = 7'h28 == _myNewVec_39_T_3[6:0] ? myVec_40 : _GEN_11473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11475 = 7'h29 == _myNewVec_39_T_3[6:0] ? myVec_41 : _GEN_11474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11476 = 7'h2a == _myNewVec_39_T_3[6:0] ? myVec_42 : _GEN_11475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11477 = 7'h2b == _myNewVec_39_T_3[6:0] ? myVec_43 : _GEN_11476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11478 = 7'h2c == _myNewVec_39_T_3[6:0] ? myVec_44 : _GEN_11477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11479 = 7'h2d == _myNewVec_39_T_3[6:0] ? myVec_45 : _GEN_11478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11480 = 7'h2e == _myNewVec_39_T_3[6:0] ? myVec_46 : _GEN_11479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11481 = 7'h2f == _myNewVec_39_T_3[6:0] ? myVec_47 : _GEN_11480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11482 = 7'h30 == _myNewVec_39_T_3[6:0] ? myVec_48 : _GEN_11481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11483 = 7'h31 == _myNewVec_39_T_3[6:0] ? myVec_49 : _GEN_11482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11484 = 7'h32 == _myNewVec_39_T_3[6:0] ? myVec_50 : _GEN_11483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11485 = 7'h33 == _myNewVec_39_T_3[6:0] ? myVec_51 : _GEN_11484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11486 = 7'h34 == _myNewVec_39_T_3[6:0] ? myVec_52 : _GEN_11485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11487 = 7'h35 == _myNewVec_39_T_3[6:0] ? myVec_53 : _GEN_11486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11488 = 7'h36 == _myNewVec_39_T_3[6:0] ? myVec_54 : _GEN_11487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11489 = 7'h37 == _myNewVec_39_T_3[6:0] ? myVec_55 : _GEN_11488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11490 = 7'h38 == _myNewVec_39_T_3[6:0] ? myVec_56 : _GEN_11489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11491 = 7'h39 == _myNewVec_39_T_3[6:0] ? myVec_57 : _GEN_11490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11492 = 7'h3a == _myNewVec_39_T_3[6:0] ? myVec_58 : _GEN_11491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11493 = 7'h3b == _myNewVec_39_T_3[6:0] ? myVec_59 : _GEN_11492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11494 = 7'h3c == _myNewVec_39_T_3[6:0] ? myVec_60 : _GEN_11493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11495 = 7'h3d == _myNewVec_39_T_3[6:0] ? myVec_61 : _GEN_11494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11496 = 7'h3e == _myNewVec_39_T_3[6:0] ? myVec_62 : _GEN_11495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11497 = 7'h3f == _myNewVec_39_T_3[6:0] ? myVec_63 : _GEN_11496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11498 = 7'h40 == _myNewVec_39_T_3[6:0] ? myVec_64 : _GEN_11497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11499 = 7'h41 == _myNewVec_39_T_3[6:0] ? myVec_65 : _GEN_11498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11500 = 7'h42 == _myNewVec_39_T_3[6:0] ? myVec_66 : _GEN_11499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11501 = 7'h43 == _myNewVec_39_T_3[6:0] ? myVec_67 : _GEN_11500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11502 = 7'h44 == _myNewVec_39_T_3[6:0] ? myVec_68 : _GEN_11501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11503 = 7'h45 == _myNewVec_39_T_3[6:0] ? myVec_69 : _GEN_11502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11504 = 7'h46 == _myNewVec_39_T_3[6:0] ? myVec_70 : _GEN_11503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11505 = 7'h47 == _myNewVec_39_T_3[6:0] ? myVec_71 : _GEN_11504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11506 = 7'h48 == _myNewVec_39_T_3[6:0] ? myVec_72 : _GEN_11505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11507 = 7'h49 == _myNewVec_39_T_3[6:0] ? myVec_73 : _GEN_11506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11508 = 7'h4a == _myNewVec_39_T_3[6:0] ? myVec_74 : _GEN_11507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11509 = 7'h4b == _myNewVec_39_T_3[6:0] ? myVec_75 : _GEN_11508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11510 = 7'h4c == _myNewVec_39_T_3[6:0] ? myVec_76 : _GEN_11509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11511 = 7'h4d == _myNewVec_39_T_3[6:0] ? myVec_77 : _GEN_11510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11512 = 7'h4e == _myNewVec_39_T_3[6:0] ? myVec_78 : _GEN_11511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11513 = 7'h4f == _myNewVec_39_T_3[6:0] ? myVec_79 : _GEN_11512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11514 = 7'h50 == _myNewVec_39_T_3[6:0] ? myVec_80 : _GEN_11513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11515 = 7'h51 == _myNewVec_39_T_3[6:0] ? myVec_81 : _GEN_11514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11516 = 7'h52 == _myNewVec_39_T_3[6:0] ? myVec_82 : _GEN_11515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11517 = 7'h53 == _myNewVec_39_T_3[6:0] ? myVec_83 : _GEN_11516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11518 = 7'h54 == _myNewVec_39_T_3[6:0] ? myVec_84 : _GEN_11517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11519 = 7'h55 == _myNewVec_39_T_3[6:0] ? myVec_85 : _GEN_11518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11520 = 7'h56 == _myNewVec_39_T_3[6:0] ? myVec_86 : _GEN_11519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11521 = 7'h57 == _myNewVec_39_T_3[6:0] ? myVec_87 : _GEN_11520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11522 = 7'h58 == _myNewVec_39_T_3[6:0] ? myVec_88 : _GEN_11521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11523 = 7'h59 == _myNewVec_39_T_3[6:0] ? myVec_89 : _GEN_11522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11524 = 7'h5a == _myNewVec_39_T_3[6:0] ? myVec_90 : _GEN_11523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11525 = 7'h5b == _myNewVec_39_T_3[6:0] ? myVec_91 : _GEN_11524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11526 = 7'h5c == _myNewVec_39_T_3[6:0] ? myVec_92 : _GEN_11525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11527 = 7'h5d == _myNewVec_39_T_3[6:0] ? myVec_93 : _GEN_11526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11528 = 7'h5e == _myNewVec_39_T_3[6:0] ? myVec_94 : _GEN_11527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11529 = 7'h5f == _myNewVec_39_T_3[6:0] ? myVec_95 : _GEN_11528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11530 = 7'h60 == _myNewVec_39_T_3[6:0] ? myVec_96 : _GEN_11529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11531 = 7'h61 == _myNewVec_39_T_3[6:0] ? myVec_97 : _GEN_11530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11532 = 7'h62 == _myNewVec_39_T_3[6:0] ? myVec_98 : _GEN_11531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11533 = 7'h63 == _myNewVec_39_T_3[6:0] ? myVec_99 : _GEN_11532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11534 = 7'h64 == _myNewVec_39_T_3[6:0] ? myVec_100 : _GEN_11533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11535 = 7'h65 == _myNewVec_39_T_3[6:0] ? myVec_101 : _GEN_11534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11536 = 7'h66 == _myNewVec_39_T_3[6:0] ? myVec_102 : _GEN_11535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11537 = 7'h67 == _myNewVec_39_T_3[6:0] ? myVec_103 : _GEN_11536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11538 = 7'h68 == _myNewVec_39_T_3[6:0] ? myVec_104 : _GEN_11537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11539 = 7'h69 == _myNewVec_39_T_3[6:0] ? myVec_105 : _GEN_11538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11540 = 7'h6a == _myNewVec_39_T_3[6:0] ? myVec_106 : _GEN_11539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11541 = 7'h6b == _myNewVec_39_T_3[6:0] ? myVec_107 : _GEN_11540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11542 = 7'h6c == _myNewVec_39_T_3[6:0] ? myVec_108 : _GEN_11541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11543 = 7'h6d == _myNewVec_39_T_3[6:0] ? myVec_109 : _GEN_11542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11544 = 7'h6e == _myNewVec_39_T_3[6:0] ? myVec_110 : _GEN_11543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11545 = 7'h6f == _myNewVec_39_T_3[6:0] ? myVec_111 : _GEN_11544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11546 = 7'h70 == _myNewVec_39_T_3[6:0] ? myVec_112 : _GEN_11545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11547 = 7'h71 == _myNewVec_39_T_3[6:0] ? myVec_113 : _GEN_11546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11548 = 7'h72 == _myNewVec_39_T_3[6:0] ? myVec_114 : _GEN_11547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11549 = 7'h73 == _myNewVec_39_T_3[6:0] ? myVec_115 : _GEN_11548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11550 = 7'h74 == _myNewVec_39_T_3[6:0] ? myVec_116 : _GEN_11549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11551 = 7'h75 == _myNewVec_39_T_3[6:0] ? myVec_117 : _GEN_11550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11552 = 7'h76 == _myNewVec_39_T_3[6:0] ? myVec_118 : _GEN_11551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11553 = 7'h77 == _myNewVec_39_T_3[6:0] ? myVec_119 : _GEN_11552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11554 = 7'h78 == _myNewVec_39_T_3[6:0] ? myVec_120 : _GEN_11553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11555 = 7'h79 == _myNewVec_39_T_3[6:0] ? myVec_121 : _GEN_11554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11556 = 7'h7a == _myNewVec_39_T_3[6:0] ? myVec_122 : _GEN_11555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11557 = 7'h7b == _myNewVec_39_T_3[6:0] ? myVec_123 : _GEN_11556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11558 = 7'h7c == _myNewVec_39_T_3[6:0] ? myVec_124 : _GEN_11557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11559 = 7'h7d == _myNewVec_39_T_3[6:0] ? myVec_125 : _GEN_11558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11560 = 7'h7e == _myNewVec_39_T_3[6:0] ? myVec_126 : _GEN_11559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_39 = 7'h7f == _myNewVec_39_T_3[6:0] ? myVec_127 : _GEN_11560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_38_T_3 = _myNewVec_127_T_1 + 16'h59; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_11563 = 7'h1 == _myNewVec_38_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11564 = 7'h2 == _myNewVec_38_T_3[6:0] ? myVec_2 : _GEN_11563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11565 = 7'h3 == _myNewVec_38_T_3[6:0] ? myVec_3 : _GEN_11564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11566 = 7'h4 == _myNewVec_38_T_3[6:0] ? myVec_4 : _GEN_11565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11567 = 7'h5 == _myNewVec_38_T_3[6:0] ? myVec_5 : _GEN_11566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11568 = 7'h6 == _myNewVec_38_T_3[6:0] ? myVec_6 : _GEN_11567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11569 = 7'h7 == _myNewVec_38_T_3[6:0] ? myVec_7 : _GEN_11568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11570 = 7'h8 == _myNewVec_38_T_3[6:0] ? myVec_8 : _GEN_11569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11571 = 7'h9 == _myNewVec_38_T_3[6:0] ? myVec_9 : _GEN_11570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11572 = 7'ha == _myNewVec_38_T_3[6:0] ? myVec_10 : _GEN_11571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11573 = 7'hb == _myNewVec_38_T_3[6:0] ? myVec_11 : _GEN_11572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11574 = 7'hc == _myNewVec_38_T_3[6:0] ? myVec_12 : _GEN_11573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11575 = 7'hd == _myNewVec_38_T_3[6:0] ? myVec_13 : _GEN_11574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11576 = 7'he == _myNewVec_38_T_3[6:0] ? myVec_14 : _GEN_11575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11577 = 7'hf == _myNewVec_38_T_3[6:0] ? myVec_15 : _GEN_11576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11578 = 7'h10 == _myNewVec_38_T_3[6:0] ? myVec_16 : _GEN_11577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11579 = 7'h11 == _myNewVec_38_T_3[6:0] ? myVec_17 : _GEN_11578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11580 = 7'h12 == _myNewVec_38_T_3[6:0] ? myVec_18 : _GEN_11579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11581 = 7'h13 == _myNewVec_38_T_3[6:0] ? myVec_19 : _GEN_11580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11582 = 7'h14 == _myNewVec_38_T_3[6:0] ? myVec_20 : _GEN_11581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11583 = 7'h15 == _myNewVec_38_T_3[6:0] ? myVec_21 : _GEN_11582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11584 = 7'h16 == _myNewVec_38_T_3[6:0] ? myVec_22 : _GEN_11583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11585 = 7'h17 == _myNewVec_38_T_3[6:0] ? myVec_23 : _GEN_11584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11586 = 7'h18 == _myNewVec_38_T_3[6:0] ? myVec_24 : _GEN_11585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11587 = 7'h19 == _myNewVec_38_T_3[6:0] ? myVec_25 : _GEN_11586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11588 = 7'h1a == _myNewVec_38_T_3[6:0] ? myVec_26 : _GEN_11587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11589 = 7'h1b == _myNewVec_38_T_3[6:0] ? myVec_27 : _GEN_11588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11590 = 7'h1c == _myNewVec_38_T_3[6:0] ? myVec_28 : _GEN_11589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11591 = 7'h1d == _myNewVec_38_T_3[6:0] ? myVec_29 : _GEN_11590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11592 = 7'h1e == _myNewVec_38_T_3[6:0] ? myVec_30 : _GEN_11591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11593 = 7'h1f == _myNewVec_38_T_3[6:0] ? myVec_31 : _GEN_11592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11594 = 7'h20 == _myNewVec_38_T_3[6:0] ? myVec_32 : _GEN_11593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11595 = 7'h21 == _myNewVec_38_T_3[6:0] ? myVec_33 : _GEN_11594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11596 = 7'h22 == _myNewVec_38_T_3[6:0] ? myVec_34 : _GEN_11595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11597 = 7'h23 == _myNewVec_38_T_3[6:0] ? myVec_35 : _GEN_11596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11598 = 7'h24 == _myNewVec_38_T_3[6:0] ? myVec_36 : _GEN_11597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11599 = 7'h25 == _myNewVec_38_T_3[6:0] ? myVec_37 : _GEN_11598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11600 = 7'h26 == _myNewVec_38_T_3[6:0] ? myVec_38 : _GEN_11599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11601 = 7'h27 == _myNewVec_38_T_3[6:0] ? myVec_39 : _GEN_11600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11602 = 7'h28 == _myNewVec_38_T_3[6:0] ? myVec_40 : _GEN_11601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11603 = 7'h29 == _myNewVec_38_T_3[6:0] ? myVec_41 : _GEN_11602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11604 = 7'h2a == _myNewVec_38_T_3[6:0] ? myVec_42 : _GEN_11603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11605 = 7'h2b == _myNewVec_38_T_3[6:0] ? myVec_43 : _GEN_11604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11606 = 7'h2c == _myNewVec_38_T_3[6:0] ? myVec_44 : _GEN_11605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11607 = 7'h2d == _myNewVec_38_T_3[6:0] ? myVec_45 : _GEN_11606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11608 = 7'h2e == _myNewVec_38_T_3[6:0] ? myVec_46 : _GEN_11607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11609 = 7'h2f == _myNewVec_38_T_3[6:0] ? myVec_47 : _GEN_11608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11610 = 7'h30 == _myNewVec_38_T_3[6:0] ? myVec_48 : _GEN_11609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11611 = 7'h31 == _myNewVec_38_T_3[6:0] ? myVec_49 : _GEN_11610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11612 = 7'h32 == _myNewVec_38_T_3[6:0] ? myVec_50 : _GEN_11611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11613 = 7'h33 == _myNewVec_38_T_3[6:0] ? myVec_51 : _GEN_11612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11614 = 7'h34 == _myNewVec_38_T_3[6:0] ? myVec_52 : _GEN_11613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11615 = 7'h35 == _myNewVec_38_T_3[6:0] ? myVec_53 : _GEN_11614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11616 = 7'h36 == _myNewVec_38_T_3[6:0] ? myVec_54 : _GEN_11615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11617 = 7'h37 == _myNewVec_38_T_3[6:0] ? myVec_55 : _GEN_11616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11618 = 7'h38 == _myNewVec_38_T_3[6:0] ? myVec_56 : _GEN_11617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11619 = 7'h39 == _myNewVec_38_T_3[6:0] ? myVec_57 : _GEN_11618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11620 = 7'h3a == _myNewVec_38_T_3[6:0] ? myVec_58 : _GEN_11619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11621 = 7'h3b == _myNewVec_38_T_3[6:0] ? myVec_59 : _GEN_11620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11622 = 7'h3c == _myNewVec_38_T_3[6:0] ? myVec_60 : _GEN_11621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11623 = 7'h3d == _myNewVec_38_T_3[6:0] ? myVec_61 : _GEN_11622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11624 = 7'h3e == _myNewVec_38_T_3[6:0] ? myVec_62 : _GEN_11623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11625 = 7'h3f == _myNewVec_38_T_3[6:0] ? myVec_63 : _GEN_11624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11626 = 7'h40 == _myNewVec_38_T_3[6:0] ? myVec_64 : _GEN_11625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11627 = 7'h41 == _myNewVec_38_T_3[6:0] ? myVec_65 : _GEN_11626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11628 = 7'h42 == _myNewVec_38_T_3[6:0] ? myVec_66 : _GEN_11627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11629 = 7'h43 == _myNewVec_38_T_3[6:0] ? myVec_67 : _GEN_11628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11630 = 7'h44 == _myNewVec_38_T_3[6:0] ? myVec_68 : _GEN_11629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11631 = 7'h45 == _myNewVec_38_T_3[6:0] ? myVec_69 : _GEN_11630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11632 = 7'h46 == _myNewVec_38_T_3[6:0] ? myVec_70 : _GEN_11631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11633 = 7'h47 == _myNewVec_38_T_3[6:0] ? myVec_71 : _GEN_11632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11634 = 7'h48 == _myNewVec_38_T_3[6:0] ? myVec_72 : _GEN_11633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11635 = 7'h49 == _myNewVec_38_T_3[6:0] ? myVec_73 : _GEN_11634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11636 = 7'h4a == _myNewVec_38_T_3[6:0] ? myVec_74 : _GEN_11635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11637 = 7'h4b == _myNewVec_38_T_3[6:0] ? myVec_75 : _GEN_11636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11638 = 7'h4c == _myNewVec_38_T_3[6:0] ? myVec_76 : _GEN_11637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11639 = 7'h4d == _myNewVec_38_T_3[6:0] ? myVec_77 : _GEN_11638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11640 = 7'h4e == _myNewVec_38_T_3[6:0] ? myVec_78 : _GEN_11639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11641 = 7'h4f == _myNewVec_38_T_3[6:0] ? myVec_79 : _GEN_11640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11642 = 7'h50 == _myNewVec_38_T_3[6:0] ? myVec_80 : _GEN_11641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11643 = 7'h51 == _myNewVec_38_T_3[6:0] ? myVec_81 : _GEN_11642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11644 = 7'h52 == _myNewVec_38_T_3[6:0] ? myVec_82 : _GEN_11643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11645 = 7'h53 == _myNewVec_38_T_3[6:0] ? myVec_83 : _GEN_11644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11646 = 7'h54 == _myNewVec_38_T_3[6:0] ? myVec_84 : _GEN_11645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11647 = 7'h55 == _myNewVec_38_T_3[6:0] ? myVec_85 : _GEN_11646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11648 = 7'h56 == _myNewVec_38_T_3[6:0] ? myVec_86 : _GEN_11647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11649 = 7'h57 == _myNewVec_38_T_3[6:0] ? myVec_87 : _GEN_11648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11650 = 7'h58 == _myNewVec_38_T_3[6:0] ? myVec_88 : _GEN_11649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11651 = 7'h59 == _myNewVec_38_T_3[6:0] ? myVec_89 : _GEN_11650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11652 = 7'h5a == _myNewVec_38_T_3[6:0] ? myVec_90 : _GEN_11651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11653 = 7'h5b == _myNewVec_38_T_3[6:0] ? myVec_91 : _GEN_11652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11654 = 7'h5c == _myNewVec_38_T_3[6:0] ? myVec_92 : _GEN_11653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11655 = 7'h5d == _myNewVec_38_T_3[6:0] ? myVec_93 : _GEN_11654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11656 = 7'h5e == _myNewVec_38_T_3[6:0] ? myVec_94 : _GEN_11655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11657 = 7'h5f == _myNewVec_38_T_3[6:0] ? myVec_95 : _GEN_11656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11658 = 7'h60 == _myNewVec_38_T_3[6:0] ? myVec_96 : _GEN_11657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11659 = 7'h61 == _myNewVec_38_T_3[6:0] ? myVec_97 : _GEN_11658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11660 = 7'h62 == _myNewVec_38_T_3[6:0] ? myVec_98 : _GEN_11659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11661 = 7'h63 == _myNewVec_38_T_3[6:0] ? myVec_99 : _GEN_11660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11662 = 7'h64 == _myNewVec_38_T_3[6:0] ? myVec_100 : _GEN_11661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11663 = 7'h65 == _myNewVec_38_T_3[6:0] ? myVec_101 : _GEN_11662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11664 = 7'h66 == _myNewVec_38_T_3[6:0] ? myVec_102 : _GEN_11663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11665 = 7'h67 == _myNewVec_38_T_3[6:0] ? myVec_103 : _GEN_11664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11666 = 7'h68 == _myNewVec_38_T_3[6:0] ? myVec_104 : _GEN_11665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11667 = 7'h69 == _myNewVec_38_T_3[6:0] ? myVec_105 : _GEN_11666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11668 = 7'h6a == _myNewVec_38_T_3[6:0] ? myVec_106 : _GEN_11667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11669 = 7'h6b == _myNewVec_38_T_3[6:0] ? myVec_107 : _GEN_11668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11670 = 7'h6c == _myNewVec_38_T_3[6:0] ? myVec_108 : _GEN_11669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11671 = 7'h6d == _myNewVec_38_T_3[6:0] ? myVec_109 : _GEN_11670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11672 = 7'h6e == _myNewVec_38_T_3[6:0] ? myVec_110 : _GEN_11671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11673 = 7'h6f == _myNewVec_38_T_3[6:0] ? myVec_111 : _GEN_11672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11674 = 7'h70 == _myNewVec_38_T_3[6:0] ? myVec_112 : _GEN_11673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11675 = 7'h71 == _myNewVec_38_T_3[6:0] ? myVec_113 : _GEN_11674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11676 = 7'h72 == _myNewVec_38_T_3[6:0] ? myVec_114 : _GEN_11675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11677 = 7'h73 == _myNewVec_38_T_3[6:0] ? myVec_115 : _GEN_11676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11678 = 7'h74 == _myNewVec_38_T_3[6:0] ? myVec_116 : _GEN_11677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11679 = 7'h75 == _myNewVec_38_T_3[6:0] ? myVec_117 : _GEN_11678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11680 = 7'h76 == _myNewVec_38_T_3[6:0] ? myVec_118 : _GEN_11679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11681 = 7'h77 == _myNewVec_38_T_3[6:0] ? myVec_119 : _GEN_11680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11682 = 7'h78 == _myNewVec_38_T_3[6:0] ? myVec_120 : _GEN_11681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11683 = 7'h79 == _myNewVec_38_T_3[6:0] ? myVec_121 : _GEN_11682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11684 = 7'h7a == _myNewVec_38_T_3[6:0] ? myVec_122 : _GEN_11683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11685 = 7'h7b == _myNewVec_38_T_3[6:0] ? myVec_123 : _GEN_11684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11686 = 7'h7c == _myNewVec_38_T_3[6:0] ? myVec_124 : _GEN_11685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11687 = 7'h7d == _myNewVec_38_T_3[6:0] ? myVec_125 : _GEN_11686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11688 = 7'h7e == _myNewVec_38_T_3[6:0] ? myVec_126 : _GEN_11687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_38 = 7'h7f == _myNewVec_38_T_3[6:0] ? myVec_127 : _GEN_11688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_37_T_3 = _myNewVec_127_T_1 + 16'h5a; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_11691 = 7'h1 == _myNewVec_37_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11692 = 7'h2 == _myNewVec_37_T_3[6:0] ? myVec_2 : _GEN_11691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11693 = 7'h3 == _myNewVec_37_T_3[6:0] ? myVec_3 : _GEN_11692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11694 = 7'h4 == _myNewVec_37_T_3[6:0] ? myVec_4 : _GEN_11693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11695 = 7'h5 == _myNewVec_37_T_3[6:0] ? myVec_5 : _GEN_11694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11696 = 7'h6 == _myNewVec_37_T_3[6:0] ? myVec_6 : _GEN_11695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11697 = 7'h7 == _myNewVec_37_T_3[6:0] ? myVec_7 : _GEN_11696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11698 = 7'h8 == _myNewVec_37_T_3[6:0] ? myVec_8 : _GEN_11697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11699 = 7'h9 == _myNewVec_37_T_3[6:0] ? myVec_9 : _GEN_11698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11700 = 7'ha == _myNewVec_37_T_3[6:0] ? myVec_10 : _GEN_11699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11701 = 7'hb == _myNewVec_37_T_3[6:0] ? myVec_11 : _GEN_11700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11702 = 7'hc == _myNewVec_37_T_3[6:0] ? myVec_12 : _GEN_11701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11703 = 7'hd == _myNewVec_37_T_3[6:0] ? myVec_13 : _GEN_11702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11704 = 7'he == _myNewVec_37_T_3[6:0] ? myVec_14 : _GEN_11703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11705 = 7'hf == _myNewVec_37_T_3[6:0] ? myVec_15 : _GEN_11704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11706 = 7'h10 == _myNewVec_37_T_3[6:0] ? myVec_16 : _GEN_11705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11707 = 7'h11 == _myNewVec_37_T_3[6:0] ? myVec_17 : _GEN_11706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11708 = 7'h12 == _myNewVec_37_T_3[6:0] ? myVec_18 : _GEN_11707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11709 = 7'h13 == _myNewVec_37_T_3[6:0] ? myVec_19 : _GEN_11708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11710 = 7'h14 == _myNewVec_37_T_3[6:0] ? myVec_20 : _GEN_11709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11711 = 7'h15 == _myNewVec_37_T_3[6:0] ? myVec_21 : _GEN_11710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11712 = 7'h16 == _myNewVec_37_T_3[6:0] ? myVec_22 : _GEN_11711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11713 = 7'h17 == _myNewVec_37_T_3[6:0] ? myVec_23 : _GEN_11712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11714 = 7'h18 == _myNewVec_37_T_3[6:0] ? myVec_24 : _GEN_11713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11715 = 7'h19 == _myNewVec_37_T_3[6:0] ? myVec_25 : _GEN_11714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11716 = 7'h1a == _myNewVec_37_T_3[6:0] ? myVec_26 : _GEN_11715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11717 = 7'h1b == _myNewVec_37_T_3[6:0] ? myVec_27 : _GEN_11716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11718 = 7'h1c == _myNewVec_37_T_3[6:0] ? myVec_28 : _GEN_11717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11719 = 7'h1d == _myNewVec_37_T_3[6:0] ? myVec_29 : _GEN_11718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11720 = 7'h1e == _myNewVec_37_T_3[6:0] ? myVec_30 : _GEN_11719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11721 = 7'h1f == _myNewVec_37_T_3[6:0] ? myVec_31 : _GEN_11720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11722 = 7'h20 == _myNewVec_37_T_3[6:0] ? myVec_32 : _GEN_11721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11723 = 7'h21 == _myNewVec_37_T_3[6:0] ? myVec_33 : _GEN_11722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11724 = 7'h22 == _myNewVec_37_T_3[6:0] ? myVec_34 : _GEN_11723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11725 = 7'h23 == _myNewVec_37_T_3[6:0] ? myVec_35 : _GEN_11724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11726 = 7'h24 == _myNewVec_37_T_3[6:0] ? myVec_36 : _GEN_11725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11727 = 7'h25 == _myNewVec_37_T_3[6:0] ? myVec_37 : _GEN_11726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11728 = 7'h26 == _myNewVec_37_T_3[6:0] ? myVec_38 : _GEN_11727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11729 = 7'h27 == _myNewVec_37_T_3[6:0] ? myVec_39 : _GEN_11728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11730 = 7'h28 == _myNewVec_37_T_3[6:0] ? myVec_40 : _GEN_11729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11731 = 7'h29 == _myNewVec_37_T_3[6:0] ? myVec_41 : _GEN_11730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11732 = 7'h2a == _myNewVec_37_T_3[6:0] ? myVec_42 : _GEN_11731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11733 = 7'h2b == _myNewVec_37_T_3[6:0] ? myVec_43 : _GEN_11732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11734 = 7'h2c == _myNewVec_37_T_3[6:0] ? myVec_44 : _GEN_11733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11735 = 7'h2d == _myNewVec_37_T_3[6:0] ? myVec_45 : _GEN_11734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11736 = 7'h2e == _myNewVec_37_T_3[6:0] ? myVec_46 : _GEN_11735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11737 = 7'h2f == _myNewVec_37_T_3[6:0] ? myVec_47 : _GEN_11736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11738 = 7'h30 == _myNewVec_37_T_3[6:0] ? myVec_48 : _GEN_11737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11739 = 7'h31 == _myNewVec_37_T_3[6:0] ? myVec_49 : _GEN_11738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11740 = 7'h32 == _myNewVec_37_T_3[6:0] ? myVec_50 : _GEN_11739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11741 = 7'h33 == _myNewVec_37_T_3[6:0] ? myVec_51 : _GEN_11740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11742 = 7'h34 == _myNewVec_37_T_3[6:0] ? myVec_52 : _GEN_11741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11743 = 7'h35 == _myNewVec_37_T_3[6:0] ? myVec_53 : _GEN_11742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11744 = 7'h36 == _myNewVec_37_T_3[6:0] ? myVec_54 : _GEN_11743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11745 = 7'h37 == _myNewVec_37_T_3[6:0] ? myVec_55 : _GEN_11744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11746 = 7'h38 == _myNewVec_37_T_3[6:0] ? myVec_56 : _GEN_11745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11747 = 7'h39 == _myNewVec_37_T_3[6:0] ? myVec_57 : _GEN_11746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11748 = 7'h3a == _myNewVec_37_T_3[6:0] ? myVec_58 : _GEN_11747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11749 = 7'h3b == _myNewVec_37_T_3[6:0] ? myVec_59 : _GEN_11748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11750 = 7'h3c == _myNewVec_37_T_3[6:0] ? myVec_60 : _GEN_11749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11751 = 7'h3d == _myNewVec_37_T_3[6:0] ? myVec_61 : _GEN_11750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11752 = 7'h3e == _myNewVec_37_T_3[6:0] ? myVec_62 : _GEN_11751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11753 = 7'h3f == _myNewVec_37_T_3[6:0] ? myVec_63 : _GEN_11752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11754 = 7'h40 == _myNewVec_37_T_3[6:0] ? myVec_64 : _GEN_11753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11755 = 7'h41 == _myNewVec_37_T_3[6:0] ? myVec_65 : _GEN_11754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11756 = 7'h42 == _myNewVec_37_T_3[6:0] ? myVec_66 : _GEN_11755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11757 = 7'h43 == _myNewVec_37_T_3[6:0] ? myVec_67 : _GEN_11756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11758 = 7'h44 == _myNewVec_37_T_3[6:0] ? myVec_68 : _GEN_11757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11759 = 7'h45 == _myNewVec_37_T_3[6:0] ? myVec_69 : _GEN_11758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11760 = 7'h46 == _myNewVec_37_T_3[6:0] ? myVec_70 : _GEN_11759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11761 = 7'h47 == _myNewVec_37_T_3[6:0] ? myVec_71 : _GEN_11760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11762 = 7'h48 == _myNewVec_37_T_3[6:0] ? myVec_72 : _GEN_11761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11763 = 7'h49 == _myNewVec_37_T_3[6:0] ? myVec_73 : _GEN_11762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11764 = 7'h4a == _myNewVec_37_T_3[6:0] ? myVec_74 : _GEN_11763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11765 = 7'h4b == _myNewVec_37_T_3[6:0] ? myVec_75 : _GEN_11764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11766 = 7'h4c == _myNewVec_37_T_3[6:0] ? myVec_76 : _GEN_11765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11767 = 7'h4d == _myNewVec_37_T_3[6:0] ? myVec_77 : _GEN_11766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11768 = 7'h4e == _myNewVec_37_T_3[6:0] ? myVec_78 : _GEN_11767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11769 = 7'h4f == _myNewVec_37_T_3[6:0] ? myVec_79 : _GEN_11768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11770 = 7'h50 == _myNewVec_37_T_3[6:0] ? myVec_80 : _GEN_11769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11771 = 7'h51 == _myNewVec_37_T_3[6:0] ? myVec_81 : _GEN_11770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11772 = 7'h52 == _myNewVec_37_T_3[6:0] ? myVec_82 : _GEN_11771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11773 = 7'h53 == _myNewVec_37_T_3[6:0] ? myVec_83 : _GEN_11772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11774 = 7'h54 == _myNewVec_37_T_3[6:0] ? myVec_84 : _GEN_11773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11775 = 7'h55 == _myNewVec_37_T_3[6:0] ? myVec_85 : _GEN_11774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11776 = 7'h56 == _myNewVec_37_T_3[6:0] ? myVec_86 : _GEN_11775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11777 = 7'h57 == _myNewVec_37_T_3[6:0] ? myVec_87 : _GEN_11776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11778 = 7'h58 == _myNewVec_37_T_3[6:0] ? myVec_88 : _GEN_11777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11779 = 7'h59 == _myNewVec_37_T_3[6:0] ? myVec_89 : _GEN_11778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11780 = 7'h5a == _myNewVec_37_T_3[6:0] ? myVec_90 : _GEN_11779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11781 = 7'h5b == _myNewVec_37_T_3[6:0] ? myVec_91 : _GEN_11780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11782 = 7'h5c == _myNewVec_37_T_3[6:0] ? myVec_92 : _GEN_11781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11783 = 7'h5d == _myNewVec_37_T_3[6:0] ? myVec_93 : _GEN_11782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11784 = 7'h5e == _myNewVec_37_T_3[6:0] ? myVec_94 : _GEN_11783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11785 = 7'h5f == _myNewVec_37_T_3[6:0] ? myVec_95 : _GEN_11784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11786 = 7'h60 == _myNewVec_37_T_3[6:0] ? myVec_96 : _GEN_11785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11787 = 7'h61 == _myNewVec_37_T_3[6:0] ? myVec_97 : _GEN_11786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11788 = 7'h62 == _myNewVec_37_T_3[6:0] ? myVec_98 : _GEN_11787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11789 = 7'h63 == _myNewVec_37_T_3[6:0] ? myVec_99 : _GEN_11788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11790 = 7'h64 == _myNewVec_37_T_3[6:0] ? myVec_100 : _GEN_11789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11791 = 7'h65 == _myNewVec_37_T_3[6:0] ? myVec_101 : _GEN_11790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11792 = 7'h66 == _myNewVec_37_T_3[6:0] ? myVec_102 : _GEN_11791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11793 = 7'h67 == _myNewVec_37_T_3[6:0] ? myVec_103 : _GEN_11792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11794 = 7'h68 == _myNewVec_37_T_3[6:0] ? myVec_104 : _GEN_11793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11795 = 7'h69 == _myNewVec_37_T_3[6:0] ? myVec_105 : _GEN_11794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11796 = 7'h6a == _myNewVec_37_T_3[6:0] ? myVec_106 : _GEN_11795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11797 = 7'h6b == _myNewVec_37_T_3[6:0] ? myVec_107 : _GEN_11796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11798 = 7'h6c == _myNewVec_37_T_3[6:0] ? myVec_108 : _GEN_11797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11799 = 7'h6d == _myNewVec_37_T_3[6:0] ? myVec_109 : _GEN_11798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11800 = 7'h6e == _myNewVec_37_T_3[6:0] ? myVec_110 : _GEN_11799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11801 = 7'h6f == _myNewVec_37_T_3[6:0] ? myVec_111 : _GEN_11800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11802 = 7'h70 == _myNewVec_37_T_3[6:0] ? myVec_112 : _GEN_11801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11803 = 7'h71 == _myNewVec_37_T_3[6:0] ? myVec_113 : _GEN_11802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11804 = 7'h72 == _myNewVec_37_T_3[6:0] ? myVec_114 : _GEN_11803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11805 = 7'h73 == _myNewVec_37_T_3[6:0] ? myVec_115 : _GEN_11804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11806 = 7'h74 == _myNewVec_37_T_3[6:0] ? myVec_116 : _GEN_11805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11807 = 7'h75 == _myNewVec_37_T_3[6:0] ? myVec_117 : _GEN_11806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11808 = 7'h76 == _myNewVec_37_T_3[6:0] ? myVec_118 : _GEN_11807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11809 = 7'h77 == _myNewVec_37_T_3[6:0] ? myVec_119 : _GEN_11808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11810 = 7'h78 == _myNewVec_37_T_3[6:0] ? myVec_120 : _GEN_11809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11811 = 7'h79 == _myNewVec_37_T_3[6:0] ? myVec_121 : _GEN_11810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11812 = 7'h7a == _myNewVec_37_T_3[6:0] ? myVec_122 : _GEN_11811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11813 = 7'h7b == _myNewVec_37_T_3[6:0] ? myVec_123 : _GEN_11812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11814 = 7'h7c == _myNewVec_37_T_3[6:0] ? myVec_124 : _GEN_11813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11815 = 7'h7d == _myNewVec_37_T_3[6:0] ? myVec_125 : _GEN_11814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11816 = 7'h7e == _myNewVec_37_T_3[6:0] ? myVec_126 : _GEN_11815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_37 = 7'h7f == _myNewVec_37_T_3[6:0] ? myVec_127 : _GEN_11816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_36_T_3 = _myNewVec_127_T_1 + 16'h5b; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_11819 = 7'h1 == _myNewVec_36_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11820 = 7'h2 == _myNewVec_36_T_3[6:0] ? myVec_2 : _GEN_11819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11821 = 7'h3 == _myNewVec_36_T_3[6:0] ? myVec_3 : _GEN_11820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11822 = 7'h4 == _myNewVec_36_T_3[6:0] ? myVec_4 : _GEN_11821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11823 = 7'h5 == _myNewVec_36_T_3[6:0] ? myVec_5 : _GEN_11822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11824 = 7'h6 == _myNewVec_36_T_3[6:0] ? myVec_6 : _GEN_11823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11825 = 7'h7 == _myNewVec_36_T_3[6:0] ? myVec_7 : _GEN_11824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11826 = 7'h8 == _myNewVec_36_T_3[6:0] ? myVec_8 : _GEN_11825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11827 = 7'h9 == _myNewVec_36_T_3[6:0] ? myVec_9 : _GEN_11826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11828 = 7'ha == _myNewVec_36_T_3[6:0] ? myVec_10 : _GEN_11827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11829 = 7'hb == _myNewVec_36_T_3[6:0] ? myVec_11 : _GEN_11828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11830 = 7'hc == _myNewVec_36_T_3[6:0] ? myVec_12 : _GEN_11829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11831 = 7'hd == _myNewVec_36_T_3[6:0] ? myVec_13 : _GEN_11830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11832 = 7'he == _myNewVec_36_T_3[6:0] ? myVec_14 : _GEN_11831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11833 = 7'hf == _myNewVec_36_T_3[6:0] ? myVec_15 : _GEN_11832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11834 = 7'h10 == _myNewVec_36_T_3[6:0] ? myVec_16 : _GEN_11833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11835 = 7'h11 == _myNewVec_36_T_3[6:0] ? myVec_17 : _GEN_11834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11836 = 7'h12 == _myNewVec_36_T_3[6:0] ? myVec_18 : _GEN_11835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11837 = 7'h13 == _myNewVec_36_T_3[6:0] ? myVec_19 : _GEN_11836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11838 = 7'h14 == _myNewVec_36_T_3[6:0] ? myVec_20 : _GEN_11837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11839 = 7'h15 == _myNewVec_36_T_3[6:0] ? myVec_21 : _GEN_11838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11840 = 7'h16 == _myNewVec_36_T_3[6:0] ? myVec_22 : _GEN_11839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11841 = 7'h17 == _myNewVec_36_T_3[6:0] ? myVec_23 : _GEN_11840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11842 = 7'h18 == _myNewVec_36_T_3[6:0] ? myVec_24 : _GEN_11841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11843 = 7'h19 == _myNewVec_36_T_3[6:0] ? myVec_25 : _GEN_11842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11844 = 7'h1a == _myNewVec_36_T_3[6:0] ? myVec_26 : _GEN_11843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11845 = 7'h1b == _myNewVec_36_T_3[6:0] ? myVec_27 : _GEN_11844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11846 = 7'h1c == _myNewVec_36_T_3[6:0] ? myVec_28 : _GEN_11845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11847 = 7'h1d == _myNewVec_36_T_3[6:0] ? myVec_29 : _GEN_11846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11848 = 7'h1e == _myNewVec_36_T_3[6:0] ? myVec_30 : _GEN_11847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11849 = 7'h1f == _myNewVec_36_T_3[6:0] ? myVec_31 : _GEN_11848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11850 = 7'h20 == _myNewVec_36_T_3[6:0] ? myVec_32 : _GEN_11849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11851 = 7'h21 == _myNewVec_36_T_3[6:0] ? myVec_33 : _GEN_11850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11852 = 7'h22 == _myNewVec_36_T_3[6:0] ? myVec_34 : _GEN_11851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11853 = 7'h23 == _myNewVec_36_T_3[6:0] ? myVec_35 : _GEN_11852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11854 = 7'h24 == _myNewVec_36_T_3[6:0] ? myVec_36 : _GEN_11853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11855 = 7'h25 == _myNewVec_36_T_3[6:0] ? myVec_37 : _GEN_11854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11856 = 7'h26 == _myNewVec_36_T_3[6:0] ? myVec_38 : _GEN_11855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11857 = 7'h27 == _myNewVec_36_T_3[6:0] ? myVec_39 : _GEN_11856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11858 = 7'h28 == _myNewVec_36_T_3[6:0] ? myVec_40 : _GEN_11857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11859 = 7'h29 == _myNewVec_36_T_3[6:0] ? myVec_41 : _GEN_11858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11860 = 7'h2a == _myNewVec_36_T_3[6:0] ? myVec_42 : _GEN_11859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11861 = 7'h2b == _myNewVec_36_T_3[6:0] ? myVec_43 : _GEN_11860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11862 = 7'h2c == _myNewVec_36_T_3[6:0] ? myVec_44 : _GEN_11861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11863 = 7'h2d == _myNewVec_36_T_3[6:0] ? myVec_45 : _GEN_11862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11864 = 7'h2e == _myNewVec_36_T_3[6:0] ? myVec_46 : _GEN_11863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11865 = 7'h2f == _myNewVec_36_T_3[6:0] ? myVec_47 : _GEN_11864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11866 = 7'h30 == _myNewVec_36_T_3[6:0] ? myVec_48 : _GEN_11865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11867 = 7'h31 == _myNewVec_36_T_3[6:0] ? myVec_49 : _GEN_11866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11868 = 7'h32 == _myNewVec_36_T_3[6:0] ? myVec_50 : _GEN_11867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11869 = 7'h33 == _myNewVec_36_T_3[6:0] ? myVec_51 : _GEN_11868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11870 = 7'h34 == _myNewVec_36_T_3[6:0] ? myVec_52 : _GEN_11869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11871 = 7'h35 == _myNewVec_36_T_3[6:0] ? myVec_53 : _GEN_11870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11872 = 7'h36 == _myNewVec_36_T_3[6:0] ? myVec_54 : _GEN_11871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11873 = 7'h37 == _myNewVec_36_T_3[6:0] ? myVec_55 : _GEN_11872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11874 = 7'h38 == _myNewVec_36_T_3[6:0] ? myVec_56 : _GEN_11873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11875 = 7'h39 == _myNewVec_36_T_3[6:0] ? myVec_57 : _GEN_11874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11876 = 7'h3a == _myNewVec_36_T_3[6:0] ? myVec_58 : _GEN_11875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11877 = 7'h3b == _myNewVec_36_T_3[6:0] ? myVec_59 : _GEN_11876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11878 = 7'h3c == _myNewVec_36_T_3[6:0] ? myVec_60 : _GEN_11877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11879 = 7'h3d == _myNewVec_36_T_3[6:0] ? myVec_61 : _GEN_11878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11880 = 7'h3e == _myNewVec_36_T_3[6:0] ? myVec_62 : _GEN_11879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11881 = 7'h3f == _myNewVec_36_T_3[6:0] ? myVec_63 : _GEN_11880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11882 = 7'h40 == _myNewVec_36_T_3[6:0] ? myVec_64 : _GEN_11881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11883 = 7'h41 == _myNewVec_36_T_3[6:0] ? myVec_65 : _GEN_11882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11884 = 7'h42 == _myNewVec_36_T_3[6:0] ? myVec_66 : _GEN_11883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11885 = 7'h43 == _myNewVec_36_T_3[6:0] ? myVec_67 : _GEN_11884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11886 = 7'h44 == _myNewVec_36_T_3[6:0] ? myVec_68 : _GEN_11885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11887 = 7'h45 == _myNewVec_36_T_3[6:0] ? myVec_69 : _GEN_11886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11888 = 7'h46 == _myNewVec_36_T_3[6:0] ? myVec_70 : _GEN_11887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11889 = 7'h47 == _myNewVec_36_T_3[6:0] ? myVec_71 : _GEN_11888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11890 = 7'h48 == _myNewVec_36_T_3[6:0] ? myVec_72 : _GEN_11889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11891 = 7'h49 == _myNewVec_36_T_3[6:0] ? myVec_73 : _GEN_11890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11892 = 7'h4a == _myNewVec_36_T_3[6:0] ? myVec_74 : _GEN_11891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11893 = 7'h4b == _myNewVec_36_T_3[6:0] ? myVec_75 : _GEN_11892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11894 = 7'h4c == _myNewVec_36_T_3[6:0] ? myVec_76 : _GEN_11893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11895 = 7'h4d == _myNewVec_36_T_3[6:0] ? myVec_77 : _GEN_11894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11896 = 7'h4e == _myNewVec_36_T_3[6:0] ? myVec_78 : _GEN_11895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11897 = 7'h4f == _myNewVec_36_T_3[6:0] ? myVec_79 : _GEN_11896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11898 = 7'h50 == _myNewVec_36_T_3[6:0] ? myVec_80 : _GEN_11897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11899 = 7'h51 == _myNewVec_36_T_3[6:0] ? myVec_81 : _GEN_11898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11900 = 7'h52 == _myNewVec_36_T_3[6:0] ? myVec_82 : _GEN_11899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11901 = 7'h53 == _myNewVec_36_T_3[6:0] ? myVec_83 : _GEN_11900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11902 = 7'h54 == _myNewVec_36_T_3[6:0] ? myVec_84 : _GEN_11901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11903 = 7'h55 == _myNewVec_36_T_3[6:0] ? myVec_85 : _GEN_11902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11904 = 7'h56 == _myNewVec_36_T_3[6:0] ? myVec_86 : _GEN_11903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11905 = 7'h57 == _myNewVec_36_T_3[6:0] ? myVec_87 : _GEN_11904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11906 = 7'h58 == _myNewVec_36_T_3[6:0] ? myVec_88 : _GEN_11905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11907 = 7'h59 == _myNewVec_36_T_3[6:0] ? myVec_89 : _GEN_11906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11908 = 7'h5a == _myNewVec_36_T_3[6:0] ? myVec_90 : _GEN_11907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11909 = 7'h5b == _myNewVec_36_T_3[6:0] ? myVec_91 : _GEN_11908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11910 = 7'h5c == _myNewVec_36_T_3[6:0] ? myVec_92 : _GEN_11909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11911 = 7'h5d == _myNewVec_36_T_3[6:0] ? myVec_93 : _GEN_11910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11912 = 7'h5e == _myNewVec_36_T_3[6:0] ? myVec_94 : _GEN_11911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11913 = 7'h5f == _myNewVec_36_T_3[6:0] ? myVec_95 : _GEN_11912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11914 = 7'h60 == _myNewVec_36_T_3[6:0] ? myVec_96 : _GEN_11913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11915 = 7'h61 == _myNewVec_36_T_3[6:0] ? myVec_97 : _GEN_11914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11916 = 7'h62 == _myNewVec_36_T_3[6:0] ? myVec_98 : _GEN_11915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11917 = 7'h63 == _myNewVec_36_T_3[6:0] ? myVec_99 : _GEN_11916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11918 = 7'h64 == _myNewVec_36_T_3[6:0] ? myVec_100 : _GEN_11917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11919 = 7'h65 == _myNewVec_36_T_3[6:0] ? myVec_101 : _GEN_11918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11920 = 7'h66 == _myNewVec_36_T_3[6:0] ? myVec_102 : _GEN_11919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11921 = 7'h67 == _myNewVec_36_T_3[6:0] ? myVec_103 : _GEN_11920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11922 = 7'h68 == _myNewVec_36_T_3[6:0] ? myVec_104 : _GEN_11921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11923 = 7'h69 == _myNewVec_36_T_3[6:0] ? myVec_105 : _GEN_11922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11924 = 7'h6a == _myNewVec_36_T_3[6:0] ? myVec_106 : _GEN_11923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11925 = 7'h6b == _myNewVec_36_T_3[6:0] ? myVec_107 : _GEN_11924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11926 = 7'h6c == _myNewVec_36_T_3[6:0] ? myVec_108 : _GEN_11925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11927 = 7'h6d == _myNewVec_36_T_3[6:0] ? myVec_109 : _GEN_11926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11928 = 7'h6e == _myNewVec_36_T_3[6:0] ? myVec_110 : _GEN_11927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11929 = 7'h6f == _myNewVec_36_T_3[6:0] ? myVec_111 : _GEN_11928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11930 = 7'h70 == _myNewVec_36_T_3[6:0] ? myVec_112 : _GEN_11929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11931 = 7'h71 == _myNewVec_36_T_3[6:0] ? myVec_113 : _GEN_11930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11932 = 7'h72 == _myNewVec_36_T_3[6:0] ? myVec_114 : _GEN_11931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11933 = 7'h73 == _myNewVec_36_T_3[6:0] ? myVec_115 : _GEN_11932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11934 = 7'h74 == _myNewVec_36_T_3[6:0] ? myVec_116 : _GEN_11933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11935 = 7'h75 == _myNewVec_36_T_3[6:0] ? myVec_117 : _GEN_11934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11936 = 7'h76 == _myNewVec_36_T_3[6:0] ? myVec_118 : _GEN_11935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11937 = 7'h77 == _myNewVec_36_T_3[6:0] ? myVec_119 : _GEN_11936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11938 = 7'h78 == _myNewVec_36_T_3[6:0] ? myVec_120 : _GEN_11937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11939 = 7'h79 == _myNewVec_36_T_3[6:0] ? myVec_121 : _GEN_11938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11940 = 7'h7a == _myNewVec_36_T_3[6:0] ? myVec_122 : _GEN_11939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11941 = 7'h7b == _myNewVec_36_T_3[6:0] ? myVec_123 : _GEN_11940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11942 = 7'h7c == _myNewVec_36_T_3[6:0] ? myVec_124 : _GEN_11941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11943 = 7'h7d == _myNewVec_36_T_3[6:0] ? myVec_125 : _GEN_11942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11944 = 7'h7e == _myNewVec_36_T_3[6:0] ? myVec_126 : _GEN_11943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_36 = 7'h7f == _myNewVec_36_T_3[6:0] ? myVec_127 : _GEN_11944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_35_T_3 = _myNewVec_127_T_1 + 16'h5c; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_11947 = 7'h1 == _myNewVec_35_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11948 = 7'h2 == _myNewVec_35_T_3[6:0] ? myVec_2 : _GEN_11947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11949 = 7'h3 == _myNewVec_35_T_3[6:0] ? myVec_3 : _GEN_11948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11950 = 7'h4 == _myNewVec_35_T_3[6:0] ? myVec_4 : _GEN_11949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11951 = 7'h5 == _myNewVec_35_T_3[6:0] ? myVec_5 : _GEN_11950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11952 = 7'h6 == _myNewVec_35_T_3[6:0] ? myVec_6 : _GEN_11951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11953 = 7'h7 == _myNewVec_35_T_3[6:0] ? myVec_7 : _GEN_11952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11954 = 7'h8 == _myNewVec_35_T_3[6:0] ? myVec_8 : _GEN_11953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11955 = 7'h9 == _myNewVec_35_T_3[6:0] ? myVec_9 : _GEN_11954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11956 = 7'ha == _myNewVec_35_T_3[6:0] ? myVec_10 : _GEN_11955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11957 = 7'hb == _myNewVec_35_T_3[6:0] ? myVec_11 : _GEN_11956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11958 = 7'hc == _myNewVec_35_T_3[6:0] ? myVec_12 : _GEN_11957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11959 = 7'hd == _myNewVec_35_T_3[6:0] ? myVec_13 : _GEN_11958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11960 = 7'he == _myNewVec_35_T_3[6:0] ? myVec_14 : _GEN_11959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11961 = 7'hf == _myNewVec_35_T_3[6:0] ? myVec_15 : _GEN_11960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11962 = 7'h10 == _myNewVec_35_T_3[6:0] ? myVec_16 : _GEN_11961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11963 = 7'h11 == _myNewVec_35_T_3[6:0] ? myVec_17 : _GEN_11962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11964 = 7'h12 == _myNewVec_35_T_3[6:0] ? myVec_18 : _GEN_11963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11965 = 7'h13 == _myNewVec_35_T_3[6:0] ? myVec_19 : _GEN_11964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11966 = 7'h14 == _myNewVec_35_T_3[6:0] ? myVec_20 : _GEN_11965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11967 = 7'h15 == _myNewVec_35_T_3[6:0] ? myVec_21 : _GEN_11966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11968 = 7'h16 == _myNewVec_35_T_3[6:0] ? myVec_22 : _GEN_11967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11969 = 7'h17 == _myNewVec_35_T_3[6:0] ? myVec_23 : _GEN_11968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11970 = 7'h18 == _myNewVec_35_T_3[6:0] ? myVec_24 : _GEN_11969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11971 = 7'h19 == _myNewVec_35_T_3[6:0] ? myVec_25 : _GEN_11970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11972 = 7'h1a == _myNewVec_35_T_3[6:0] ? myVec_26 : _GEN_11971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11973 = 7'h1b == _myNewVec_35_T_3[6:0] ? myVec_27 : _GEN_11972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11974 = 7'h1c == _myNewVec_35_T_3[6:0] ? myVec_28 : _GEN_11973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11975 = 7'h1d == _myNewVec_35_T_3[6:0] ? myVec_29 : _GEN_11974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11976 = 7'h1e == _myNewVec_35_T_3[6:0] ? myVec_30 : _GEN_11975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11977 = 7'h1f == _myNewVec_35_T_3[6:0] ? myVec_31 : _GEN_11976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11978 = 7'h20 == _myNewVec_35_T_3[6:0] ? myVec_32 : _GEN_11977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11979 = 7'h21 == _myNewVec_35_T_3[6:0] ? myVec_33 : _GEN_11978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11980 = 7'h22 == _myNewVec_35_T_3[6:0] ? myVec_34 : _GEN_11979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11981 = 7'h23 == _myNewVec_35_T_3[6:0] ? myVec_35 : _GEN_11980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11982 = 7'h24 == _myNewVec_35_T_3[6:0] ? myVec_36 : _GEN_11981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11983 = 7'h25 == _myNewVec_35_T_3[6:0] ? myVec_37 : _GEN_11982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11984 = 7'h26 == _myNewVec_35_T_3[6:0] ? myVec_38 : _GEN_11983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11985 = 7'h27 == _myNewVec_35_T_3[6:0] ? myVec_39 : _GEN_11984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11986 = 7'h28 == _myNewVec_35_T_3[6:0] ? myVec_40 : _GEN_11985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11987 = 7'h29 == _myNewVec_35_T_3[6:0] ? myVec_41 : _GEN_11986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11988 = 7'h2a == _myNewVec_35_T_3[6:0] ? myVec_42 : _GEN_11987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11989 = 7'h2b == _myNewVec_35_T_3[6:0] ? myVec_43 : _GEN_11988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11990 = 7'h2c == _myNewVec_35_T_3[6:0] ? myVec_44 : _GEN_11989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11991 = 7'h2d == _myNewVec_35_T_3[6:0] ? myVec_45 : _GEN_11990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11992 = 7'h2e == _myNewVec_35_T_3[6:0] ? myVec_46 : _GEN_11991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11993 = 7'h2f == _myNewVec_35_T_3[6:0] ? myVec_47 : _GEN_11992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11994 = 7'h30 == _myNewVec_35_T_3[6:0] ? myVec_48 : _GEN_11993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11995 = 7'h31 == _myNewVec_35_T_3[6:0] ? myVec_49 : _GEN_11994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11996 = 7'h32 == _myNewVec_35_T_3[6:0] ? myVec_50 : _GEN_11995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11997 = 7'h33 == _myNewVec_35_T_3[6:0] ? myVec_51 : _GEN_11996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11998 = 7'h34 == _myNewVec_35_T_3[6:0] ? myVec_52 : _GEN_11997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_11999 = 7'h35 == _myNewVec_35_T_3[6:0] ? myVec_53 : _GEN_11998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12000 = 7'h36 == _myNewVec_35_T_3[6:0] ? myVec_54 : _GEN_11999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12001 = 7'h37 == _myNewVec_35_T_3[6:0] ? myVec_55 : _GEN_12000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12002 = 7'h38 == _myNewVec_35_T_3[6:0] ? myVec_56 : _GEN_12001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12003 = 7'h39 == _myNewVec_35_T_3[6:0] ? myVec_57 : _GEN_12002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12004 = 7'h3a == _myNewVec_35_T_3[6:0] ? myVec_58 : _GEN_12003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12005 = 7'h3b == _myNewVec_35_T_3[6:0] ? myVec_59 : _GEN_12004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12006 = 7'h3c == _myNewVec_35_T_3[6:0] ? myVec_60 : _GEN_12005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12007 = 7'h3d == _myNewVec_35_T_3[6:0] ? myVec_61 : _GEN_12006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12008 = 7'h3e == _myNewVec_35_T_3[6:0] ? myVec_62 : _GEN_12007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12009 = 7'h3f == _myNewVec_35_T_3[6:0] ? myVec_63 : _GEN_12008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12010 = 7'h40 == _myNewVec_35_T_3[6:0] ? myVec_64 : _GEN_12009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12011 = 7'h41 == _myNewVec_35_T_3[6:0] ? myVec_65 : _GEN_12010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12012 = 7'h42 == _myNewVec_35_T_3[6:0] ? myVec_66 : _GEN_12011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12013 = 7'h43 == _myNewVec_35_T_3[6:0] ? myVec_67 : _GEN_12012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12014 = 7'h44 == _myNewVec_35_T_3[6:0] ? myVec_68 : _GEN_12013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12015 = 7'h45 == _myNewVec_35_T_3[6:0] ? myVec_69 : _GEN_12014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12016 = 7'h46 == _myNewVec_35_T_3[6:0] ? myVec_70 : _GEN_12015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12017 = 7'h47 == _myNewVec_35_T_3[6:0] ? myVec_71 : _GEN_12016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12018 = 7'h48 == _myNewVec_35_T_3[6:0] ? myVec_72 : _GEN_12017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12019 = 7'h49 == _myNewVec_35_T_3[6:0] ? myVec_73 : _GEN_12018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12020 = 7'h4a == _myNewVec_35_T_3[6:0] ? myVec_74 : _GEN_12019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12021 = 7'h4b == _myNewVec_35_T_3[6:0] ? myVec_75 : _GEN_12020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12022 = 7'h4c == _myNewVec_35_T_3[6:0] ? myVec_76 : _GEN_12021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12023 = 7'h4d == _myNewVec_35_T_3[6:0] ? myVec_77 : _GEN_12022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12024 = 7'h4e == _myNewVec_35_T_3[6:0] ? myVec_78 : _GEN_12023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12025 = 7'h4f == _myNewVec_35_T_3[6:0] ? myVec_79 : _GEN_12024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12026 = 7'h50 == _myNewVec_35_T_3[6:0] ? myVec_80 : _GEN_12025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12027 = 7'h51 == _myNewVec_35_T_3[6:0] ? myVec_81 : _GEN_12026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12028 = 7'h52 == _myNewVec_35_T_3[6:0] ? myVec_82 : _GEN_12027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12029 = 7'h53 == _myNewVec_35_T_3[6:0] ? myVec_83 : _GEN_12028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12030 = 7'h54 == _myNewVec_35_T_3[6:0] ? myVec_84 : _GEN_12029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12031 = 7'h55 == _myNewVec_35_T_3[6:0] ? myVec_85 : _GEN_12030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12032 = 7'h56 == _myNewVec_35_T_3[6:0] ? myVec_86 : _GEN_12031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12033 = 7'h57 == _myNewVec_35_T_3[6:0] ? myVec_87 : _GEN_12032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12034 = 7'h58 == _myNewVec_35_T_3[6:0] ? myVec_88 : _GEN_12033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12035 = 7'h59 == _myNewVec_35_T_3[6:0] ? myVec_89 : _GEN_12034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12036 = 7'h5a == _myNewVec_35_T_3[6:0] ? myVec_90 : _GEN_12035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12037 = 7'h5b == _myNewVec_35_T_3[6:0] ? myVec_91 : _GEN_12036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12038 = 7'h5c == _myNewVec_35_T_3[6:0] ? myVec_92 : _GEN_12037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12039 = 7'h5d == _myNewVec_35_T_3[6:0] ? myVec_93 : _GEN_12038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12040 = 7'h5e == _myNewVec_35_T_3[6:0] ? myVec_94 : _GEN_12039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12041 = 7'h5f == _myNewVec_35_T_3[6:0] ? myVec_95 : _GEN_12040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12042 = 7'h60 == _myNewVec_35_T_3[6:0] ? myVec_96 : _GEN_12041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12043 = 7'h61 == _myNewVec_35_T_3[6:0] ? myVec_97 : _GEN_12042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12044 = 7'h62 == _myNewVec_35_T_3[6:0] ? myVec_98 : _GEN_12043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12045 = 7'h63 == _myNewVec_35_T_3[6:0] ? myVec_99 : _GEN_12044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12046 = 7'h64 == _myNewVec_35_T_3[6:0] ? myVec_100 : _GEN_12045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12047 = 7'h65 == _myNewVec_35_T_3[6:0] ? myVec_101 : _GEN_12046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12048 = 7'h66 == _myNewVec_35_T_3[6:0] ? myVec_102 : _GEN_12047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12049 = 7'h67 == _myNewVec_35_T_3[6:0] ? myVec_103 : _GEN_12048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12050 = 7'h68 == _myNewVec_35_T_3[6:0] ? myVec_104 : _GEN_12049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12051 = 7'h69 == _myNewVec_35_T_3[6:0] ? myVec_105 : _GEN_12050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12052 = 7'h6a == _myNewVec_35_T_3[6:0] ? myVec_106 : _GEN_12051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12053 = 7'h6b == _myNewVec_35_T_3[6:0] ? myVec_107 : _GEN_12052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12054 = 7'h6c == _myNewVec_35_T_3[6:0] ? myVec_108 : _GEN_12053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12055 = 7'h6d == _myNewVec_35_T_3[6:0] ? myVec_109 : _GEN_12054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12056 = 7'h6e == _myNewVec_35_T_3[6:0] ? myVec_110 : _GEN_12055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12057 = 7'h6f == _myNewVec_35_T_3[6:0] ? myVec_111 : _GEN_12056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12058 = 7'h70 == _myNewVec_35_T_3[6:0] ? myVec_112 : _GEN_12057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12059 = 7'h71 == _myNewVec_35_T_3[6:0] ? myVec_113 : _GEN_12058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12060 = 7'h72 == _myNewVec_35_T_3[6:0] ? myVec_114 : _GEN_12059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12061 = 7'h73 == _myNewVec_35_T_3[6:0] ? myVec_115 : _GEN_12060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12062 = 7'h74 == _myNewVec_35_T_3[6:0] ? myVec_116 : _GEN_12061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12063 = 7'h75 == _myNewVec_35_T_3[6:0] ? myVec_117 : _GEN_12062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12064 = 7'h76 == _myNewVec_35_T_3[6:0] ? myVec_118 : _GEN_12063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12065 = 7'h77 == _myNewVec_35_T_3[6:0] ? myVec_119 : _GEN_12064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12066 = 7'h78 == _myNewVec_35_T_3[6:0] ? myVec_120 : _GEN_12065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12067 = 7'h79 == _myNewVec_35_T_3[6:0] ? myVec_121 : _GEN_12066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12068 = 7'h7a == _myNewVec_35_T_3[6:0] ? myVec_122 : _GEN_12067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12069 = 7'h7b == _myNewVec_35_T_3[6:0] ? myVec_123 : _GEN_12068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12070 = 7'h7c == _myNewVec_35_T_3[6:0] ? myVec_124 : _GEN_12069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12071 = 7'h7d == _myNewVec_35_T_3[6:0] ? myVec_125 : _GEN_12070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12072 = 7'h7e == _myNewVec_35_T_3[6:0] ? myVec_126 : _GEN_12071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_35 = 7'h7f == _myNewVec_35_T_3[6:0] ? myVec_127 : _GEN_12072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_34_T_3 = _myNewVec_127_T_1 + 16'h5d; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_12075 = 7'h1 == _myNewVec_34_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12076 = 7'h2 == _myNewVec_34_T_3[6:0] ? myVec_2 : _GEN_12075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12077 = 7'h3 == _myNewVec_34_T_3[6:0] ? myVec_3 : _GEN_12076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12078 = 7'h4 == _myNewVec_34_T_3[6:0] ? myVec_4 : _GEN_12077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12079 = 7'h5 == _myNewVec_34_T_3[6:0] ? myVec_5 : _GEN_12078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12080 = 7'h6 == _myNewVec_34_T_3[6:0] ? myVec_6 : _GEN_12079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12081 = 7'h7 == _myNewVec_34_T_3[6:0] ? myVec_7 : _GEN_12080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12082 = 7'h8 == _myNewVec_34_T_3[6:0] ? myVec_8 : _GEN_12081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12083 = 7'h9 == _myNewVec_34_T_3[6:0] ? myVec_9 : _GEN_12082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12084 = 7'ha == _myNewVec_34_T_3[6:0] ? myVec_10 : _GEN_12083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12085 = 7'hb == _myNewVec_34_T_3[6:0] ? myVec_11 : _GEN_12084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12086 = 7'hc == _myNewVec_34_T_3[6:0] ? myVec_12 : _GEN_12085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12087 = 7'hd == _myNewVec_34_T_3[6:0] ? myVec_13 : _GEN_12086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12088 = 7'he == _myNewVec_34_T_3[6:0] ? myVec_14 : _GEN_12087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12089 = 7'hf == _myNewVec_34_T_3[6:0] ? myVec_15 : _GEN_12088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12090 = 7'h10 == _myNewVec_34_T_3[6:0] ? myVec_16 : _GEN_12089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12091 = 7'h11 == _myNewVec_34_T_3[6:0] ? myVec_17 : _GEN_12090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12092 = 7'h12 == _myNewVec_34_T_3[6:0] ? myVec_18 : _GEN_12091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12093 = 7'h13 == _myNewVec_34_T_3[6:0] ? myVec_19 : _GEN_12092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12094 = 7'h14 == _myNewVec_34_T_3[6:0] ? myVec_20 : _GEN_12093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12095 = 7'h15 == _myNewVec_34_T_3[6:0] ? myVec_21 : _GEN_12094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12096 = 7'h16 == _myNewVec_34_T_3[6:0] ? myVec_22 : _GEN_12095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12097 = 7'h17 == _myNewVec_34_T_3[6:0] ? myVec_23 : _GEN_12096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12098 = 7'h18 == _myNewVec_34_T_3[6:0] ? myVec_24 : _GEN_12097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12099 = 7'h19 == _myNewVec_34_T_3[6:0] ? myVec_25 : _GEN_12098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12100 = 7'h1a == _myNewVec_34_T_3[6:0] ? myVec_26 : _GEN_12099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12101 = 7'h1b == _myNewVec_34_T_3[6:0] ? myVec_27 : _GEN_12100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12102 = 7'h1c == _myNewVec_34_T_3[6:0] ? myVec_28 : _GEN_12101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12103 = 7'h1d == _myNewVec_34_T_3[6:0] ? myVec_29 : _GEN_12102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12104 = 7'h1e == _myNewVec_34_T_3[6:0] ? myVec_30 : _GEN_12103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12105 = 7'h1f == _myNewVec_34_T_3[6:0] ? myVec_31 : _GEN_12104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12106 = 7'h20 == _myNewVec_34_T_3[6:0] ? myVec_32 : _GEN_12105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12107 = 7'h21 == _myNewVec_34_T_3[6:0] ? myVec_33 : _GEN_12106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12108 = 7'h22 == _myNewVec_34_T_3[6:0] ? myVec_34 : _GEN_12107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12109 = 7'h23 == _myNewVec_34_T_3[6:0] ? myVec_35 : _GEN_12108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12110 = 7'h24 == _myNewVec_34_T_3[6:0] ? myVec_36 : _GEN_12109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12111 = 7'h25 == _myNewVec_34_T_3[6:0] ? myVec_37 : _GEN_12110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12112 = 7'h26 == _myNewVec_34_T_3[6:0] ? myVec_38 : _GEN_12111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12113 = 7'h27 == _myNewVec_34_T_3[6:0] ? myVec_39 : _GEN_12112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12114 = 7'h28 == _myNewVec_34_T_3[6:0] ? myVec_40 : _GEN_12113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12115 = 7'h29 == _myNewVec_34_T_3[6:0] ? myVec_41 : _GEN_12114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12116 = 7'h2a == _myNewVec_34_T_3[6:0] ? myVec_42 : _GEN_12115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12117 = 7'h2b == _myNewVec_34_T_3[6:0] ? myVec_43 : _GEN_12116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12118 = 7'h2c == _myNewVec_34_T_3[6:0] ? myVec_44 : _GEN_12117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12119 = 7'h2d == _myNewVec_34_T_3[6:0] ? myVec_45 : _GEN_12118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12120 = 7'h2e == _myNewVec_34_T_3[6:0] ? myVec_46 : _GEN_12119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12121 = 7'h2f == _myNewVec_34_T_3[6:0] ? myVec_47 : _GEN_12120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12122 = 7'h30 == _myNewVec_34_T_3[6:0] ? myVec_48 : _GEN_12121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12123 = 7'h31 == _myNewVec_34_T_3[6:0] ? myVec_49 : _GEN_12122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12124 = 7'h32 == _myNewVec_34_T_3[6:0] ? myVec_50 : _GEN_12123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12125 = 7'h33 == _myNewVec_34_T_3[6:0] ? myVec_51 : _GEN_12124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12126 = 7'h34 == _myNewVec_34_T_3[6:0] ? myVec_52 : _GEN_12125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12127 = 7'h35 == _myNewVec_34_T_3[6:0] ? myVec_53 : _GEN_12126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12128 = 7'h36 == _myNewVec_34_T_3[6:0] ? myVec_54 : _GEN_12127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12129 = 7'h37 == _myNewVec_34_T_3[6:0] ? myVec_55 : _GEN_12128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12130 = 7'h38 == _myNewVec_34_T_3[6:0] ? myVec_56 : _GEN_12129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12131 = 7'h39 == _myNewVec_34_T_3[6:0] ? myVec_57 : _GEN_12130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12132 = 7'h3a == _myNewVec_34_T_3[6:0] ? myVec_58 : _GEN_12131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12133 = 7'h3b == _myNewVec_34_T_3[6:0] ? myVec_59 : _GEN_12132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12134 = 7'h3c == _myNewVec_34_T_3[6:0] ? myVec_60 : _GEN_12133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12135 = 7'h3d == _myNewVec_34_T_3[6:0] ? myVec_61 : _GEN_12134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12136 = 7'h3e == _myNewVec_34_T_3[6:0] ? myVec_62 : _GEN_12135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12137 = 7'h3f == _myNewVec_34_T_3[6:0] ? myVec_63 : _GEN_12136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12138 = 7'h40 == _myNewVec_34_T_3[6:0] ? myVec_64 : _GEN_12137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12139 = 7'h41 == _myNewVec_34_T_3[6:0] ? myVec_65 : _GEN_12138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12140 = 7'h42 == _myNewVec_34_T_3[6:0] ? myVec_66 : _GEN_12139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12141 = 7'h43 == _myNewVec_34_T_3[6:0] ? myVec_67 : _GEN_12140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12142 = 7'h44 == _myNewVec_34_T_3[6:0] ? myVec_68 : _GEN_12141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12143 = 7'h45 == _myNewVec_34_T_3[6:0] ? myVec_69 : _GEN_12142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12144 = 7'h46 == _myNewVec_34_T_3[6:0] ? myVec_70 : _GEN_12143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12145 = 7'h47 == _myNewVec_34_T_3[6:0] ? myVec_71 : _GEN_12144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12146 = 7'h48 == _myNewVec_34_T_3[6:0] ? myVec_72 : _GEN_12145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12147 = 7'h49 == _myNewVec_34_T_3[6:0] ? myVec_73 : _GEN_12146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12148 = 7'h4a == _myNewVec_34_T_3[6:0] ? myVec_74 : _GEN_12147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12149 = 7'h4b == _myNewVec_34_T_3[6:0] ? myVec_75 : _GEN_12148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12150 = 7'h4c == _myNewVec_34_T_3[6:0] ? myVec_76 : _GEN_12149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12151 = 7'h4d == _myNewVec_34_T_3[6:0] ? myVec_77 : _GEN_12150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12152 = 7'h4e == _myNewVec_34_T_3[6:0] ? myVec_78 : _GEN_12151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12153 = 7'h4f == _myNewVec_34_T_3[6:0] ? myVec_79 : _GEN_12152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12154 = 7'h50 == _myNewVec_34_T_3[6:0] ? myVec_80 : _GEN_12153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12155 = 7'h51 == _myNewVec_34_T_3[6:0] ? myVec_81 : _GEN_12154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12156 = 7'h52 == _myNewVec_34_T_3[6:0] ? myVec_82 : _GEN_12155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12157 = 7'h53 == _myNewVec_34_T_3[6:0] ? myVec_83 : _GEN_12156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12158 = 7'h54 == _myNewVec_34_T_3[6:0] ? myVec_84 : _GEN_12157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12159 = 7'h55 == _myNewVec_34_T_3[6:0] ? myVec_85 : _GEN_12158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12160 = 7'h56 == _myNewVec_34_T_3[6:0] ? myVec_86 : _GEN_12159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12161 = 7'h57 == _myNewVec_34_T_3[6:0] ? myVec_87 : _GEN_12160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12162 = 7'h58 == _myNewVec_34_T_3[6:0] ? myVec_88 : _GEN_12161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12163 = 7'h59 == _myNewVec_34_T_3[6:0] ? myVec_89 : _GEN_12162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12164 = 7'h5a == _myNewVec_34_T_3[6:0] ? myVec_90 : _GEN_12163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12165 = 7'h5b == _myNewVec_34_T_3[6:0] ? myVec_91 : _GEN_12164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12166 = 7'h5c == _myNewVec_34_T_3[6:0] ? myVec_92 : _GEN_12165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12167 = 7'h5d == _myNewVec_34_T_3[6:0] ? myVec_93 : _GEN_12166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12168 = 7'h5e == _myNewVec_34_T_3[6:0] ? myVec_94 : _GEN_12167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12169 = 7'h5f == _myNewVec_34_T_3[6:0] ? myVec_95 : _GEN_12168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12170 = 7'h60 == _myNewVec_34_T_3[6:0] ? myVec_96 : _GEN_12169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12171 = 7'h61 == _myNewVec_34_T_3[6:0] ? myVec_97 : _GEN_12170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12172 = 7'h62 == _myNewVec_34_T_3[6:0] ? myVec_98 : _GEN_12171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12173 = 7'h63 == _myNewVec_34_T_3[6:0] ? myVec_99 : _GEN_12172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12174 = 7'h64 == _myNewVec_34_T_3[6:0] ? myVec_100 : _GEN_12173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12175 = 7'h65 == _myNewVec_34_T_3[6:0] ? myVec_101 : _GEN_12174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12176 = 7'h66 == _myNewVec_34_T_3[6:0] ? myVec_102 : _GEN_12175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12177 = 7'h67 == _myNewVec_34_T_3[6:0] ? myVec_103 : _GEN_12176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12178 = 7'h68 == _myNewVec_34_T_3[6:0] ? myVec_104 : _GEN_12177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12179 = 7'h69 == _myNewVec_34_T_3[6:0] ? myVec_105 : _GEN_12178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12180 = 7'h6a == _myNewVec_34_T_3[6:0] ? myVec_106 : _GEN_12179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12181 = 7'h6b == _myNewVec_34_T_3[6:0] ? myVec_107 : _GEN_12180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12182 = 7'h6c == _myNewVec_34_T_3[6:0] ? myVec_108 : _GEN_12181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12183 = 7'h6d == _myNewVec_34_T_3[6:0] ? myVec_109 : _GEN_12182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12184 = 7'h6e == _myNewVec_34_T_3[6:0] ? myVec_110 : _GEN_12183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12185 = 7'h6f == _myNewVec_34_T_3[6:0] ? myVec_111 : _GEN_12184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12186 = 7'h70 == _myNewVec_34_T_3[6:0] ? myVec_112 : _GEN_12185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12187 = 7'h71 == _myNewVec_34_T_3[6:0] ? myVec_113 : _GEN_12186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12188 = 7'h72 == _myNewVec_34_T_3[6:0] ? myVec_114 : _GEN_12187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12189 = 7'h73 == _myNewVec_34_T_3[6:0] ? myVec_115 : _GEN_12188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12190 = 7'h74 == _myNewVec_34_T_3[6:0] ? myVec_116 : _GEN_12189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12191 = 7'h75 == _myNewVec_34_T_3[6:0] ? myVec_117 : _GEN_12190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12192 = 7'h76 == _myNewVec_34_T_3[6:0] ? myVec_118 : _GEN_12191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12193 = 7'h77 == _myNewVec_34_T_3[6:0] ? myVec_119 : _GEN_12192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12194 = 7'h78 == _myNewVec_34_T_3[6:0] ? myVec_120 : _GEN_12193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12195 = 7'h79 == _myNewVec_34_T_3[6:0] ? myVec_121 : _GEN_12194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12196 = 7'h7a == _myNewVec_34_T_3[6:0] ? myVec_122 : _GEN_12195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12197 = 7'h7b == _myNewVec_34_T_3[6:0] ? myVec_123 : _GEN_12196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12198 = 7'h7c == _myNewVec_34_T_3[6:0] ? myVec_124 : _GEN_12197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12199 = 7'h7d == _myNewVec_34_T_3[6:0] ? myVec_125 : _GEN_12198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12200 = 7'h7e == _myNewVec_34_T_3[6:0] ? myVec_126 : _GEN_12199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_34 = 7'h7f == _myNewVec_34_T_3[6:0] ? myVec_127 : _GEN_12200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_33_T_3 = _myNewVec_127_T_1 + 16'h5e; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_12203 = 7'h1 == _myNewVec_33_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12204 = 7'h2 == _myNewVec_33_T_3[6:0] ? myVec_2 : _GEN_12203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12205 = 7'h3 == _myNewVec_33_T_3[6:0] ? myVec_3 : _GEN_12204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12206 = 7'h4 == _myNewVec_33_T_3[6:0] ? myVec_4 : _GEN_12205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12207 = 7'h5 == _myNewVec_33_T_3[6:0] ? myVec_5 : _GEN_12206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12208 = 7'h6 == _myNewVec_33_T_3[6:0] ? myVec_6 : _GEN_12207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12209 = 7'h7 == _myNewVec_33_T_3[6:0] ? myVec_7 : _GEN_12208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12210 = 7'h8 == _myNewVec_33_T_3[6:0] ? myVec_8 : _GEN_12209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12211 = 7'h9 == _myNewVec_33_T_3[6:0] ? myVec_9 : _GEN_12210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12212 = 7'ha == _myNewVec_33_T_3[6:0] ? myVec_10 : _GEN_12211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12213 = 7'hb == _myNewVec_33_T_3[6:0] ? myVec_11 : _GEN_12212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12214 = 7'hc == _myNewVec_33_T_3[6:0] ? myVec_12 : _GEN_12213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12215 = 7'hd == _myNewVec_33_T_3[6:0] ? myVec_13 : _GEN_12214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12216 = 7'he == _myNewVec_33_T_3[6:0] ? myVec_14 : _GEN_12215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12217 = 7'hf == _myNewVec_33_T_3[6:0] ? myVec_15 : _GEN_12216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12218 = 7'h10 == _myNewVec_33_T_3[6:0] ? myVec_16 : _GEN_12217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12219 = 7'h11 == _myNewVec_33_T_3[6:0] ? myVec_17 : _GEN_12218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12220 = 7'h12 == _myNewVec_33_T_3[6:0] ? myVec_18 : _GEN_12219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12221 = 7'h13 == _myNewVec_33_T_3[6:0] ? myVec_19 : _GEN_12220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12222 = 7'h14 == _myNewVec_33_T_3[6:0] ? myVec_20 : _GEN_12221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12223 = 7'h15 == _myNewVec_33_T_3[6:0] ? myVec_21 : _GEN_12222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12224 = 7'h16 == _myNewVec_33_T_3[6:0] ? myVec_22 : _GEN_12223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12225 = 7'h17 == _myNewVec_33_T_3[6:0] ? myVec_23 : _GEN_12224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12226 = 7'h18 == _myNewVec_33_T_3[6:0] ? myVec_24 : _GEN_12225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12227 = 7'h19 == _myNewVec_33_T_3[6:0] ? myVec_25 : _GEN_12226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12228 = 7'h1a == _myNewVec_33_T_3[6:0] ? myVec_26 : _GEN_12227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12229 = 7'h1b == _myNewVec_33_T_3[6:0] ? myVec_27 : _GEN_12228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12230 = 7'h1c == _myNewVec_33_T_3[6:0] ? myVec_28 : _GEN_12229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12231 = 7'h1d == _myNewVec_33_T_3[6:0] ? myVec_29 : _GEN_12230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12232 = 7'h1e == _myNewVec_33_T_3[6:0] ? myVec_30 : _GEN_12231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12233 = 7'h1f == _myNewVec_33_T_3[6:0] ? myVec_31 : _GEN_12232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12234 = 7'h20 == _myNewVec_33_T_3[6:0] ? myVec_32 : _GEN_12233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12235 = 7'h21 == _myNewVec_33_T_3[6:0] ? myVec_33 : _GEN_12234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12236 = 7'h22 == _myNewVec_33_T_3[6:0] ? myVec_34 : _GEN_12235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12237 = 7'h23 == _myNewVec_33_T_3[6:0] ? myVec_35 : _GEN_12236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12238 = 7'h24 == _myNewVec_33_T_3[6:0] ? myVec_36 : _GEN_12237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12239 = 7'h25 == _myNewVec_33_T_3[6:0] ? myVec_37 : _GEN_12238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12240 = 7'h26 == _myNewVec_33_T_3[6:0] ? myVec_38 : _GEN_12239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12241 = 7'h27 == _myNewVec_33_T_3[6:0] ? myVec_39 : _GEN_12240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12242 = 7'h28 == _myNewVec_33_T_3[6:0] ? myVec_40 : _GEN_12241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12243 = 7'h29 == _myNewVec_33_T_3[6:0] ? myVec_41 : _GEN_12242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12244 = 7'h2a == _myNewVec_33_T_3[6:0] ? myVec_42 : _GEN_12243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12245 = 7'h2b == _myNewVec_33_T_3[6:0] ? myVec_43 : _GEN_12244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12246 = 7'h2c == _myNewVec_33_T_3[6:0] ? myVec_44 : _GEN_12245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12247 = 7'h2d == _myNewVec_33_T_3[6:0] ? myVec_45 : _GEN_12246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12248 = 7'h2e == _myNewVec_33_T_3[6:0] ? myVec_46 : _GEN_12247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12249 = 7'h2f == _myNewVec_33_T_3[6:0] ? myVec_47 : _GEN_12248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12250 = 7'h30 == _myNewVec_33_T_3[6:0] ? myVec_48 : _GEN_12249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12251 = 7'h31 == _myNewVec_33_T_3[6:0] ? myVec_49 : _GEN_12250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12252 = 7'h32 == _myNewVec_33_T_3[6:0] ? myVec_50 : _GEN_12251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12253 = 7'h33 == _myNewVec_33_T_3[6:0] ? myVec_51 : _GEN_12252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12254 = 7'h34 == _myNewVec_33_T_3[6:0] ? myVec_52 : _GEN_12253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12255 = 7'h35 == _myNewVec_33_T_3[6:0] ? myVec_53 : _GEN_12254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12256 = 7'h36 == _myNewVec_33_T_3[6:0] ? myVec_54 : _GEN_12255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12257 = 7'h37 == _myNewVec_33_T_3[6:0] ? myVec_55 : _GEN_12256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12258 = 7'h38 == _myNewVec_33_T_3[6:0] ? myVec_56 : _GEN_12257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12259 = 7'h39 == _myNewVec_33_T_3[6:0] ? myVec_57 : _GEN_12258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12260 = 7'h3a == _myNewVec_33_T_3[6:0] ? myVec_58 : _GEN_12259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12261 = 7'h3b == _myNewVec_33_T_3[6:0] ? myVec_59 : _GEN_12260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12262 = 7'h3c == _myNewVec_33_T_3[6:0] ? myVec_60 : _GEN_12261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12263 = 7'h3d == _myNewVec_33_T_3[6:0] ? myVec_61 : _GEN_12262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12264 = 7'h3e == _myNewVec_33_T_3[6:0] ? myVec_62 : _GEN_12263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12265 = 7'h3f == _myNewVec_33_T_3[6:0] ? myVec_63 : _GEN_12264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12266 = 7'h40 == _myNewVec_33_T_3[6:0] ? myVec_64 : _GEN_12265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12267 = 7'h41 == _myNewVec_33_T_3[6:0] ? myVec_65 : _GEN_12266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12268 = 7'h42 == _myNewVec_33_T_3[6:0] ? myVec_66 : _GEN_12267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12269 = 7'h43 == _myNewVec_33_T_3[6:0] ? myVec_67 : _GEN_12268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12270 = 7'h44 == _myNewVec_33_T_3[6:0] ? myVec_68 : _GEN_12269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12271 = 7'h45 == _myNewVec_33_T_3[6:0] ? myVec_69 : _GEN_12270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12272 = 7'h46 == _myNewVec_33_T_3[6:0] ? myVec_70 : _GEN_12271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12273 = 7'h47 == _myNewVec_33_T_3[6:0] ? myVec_71 : _GEN_12272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12274 = 7'h48 == _myNewVec_33_T_3[6:0] ? myVec_72 : _GEN_12273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12275 = 7'h49 == _myNewVec_33_T_3[6:0] ? myVec_73 : _GEN_12274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12276 = 7'h4a == _myNewVec_33_T_3[6:0] ? myVec_74 : _GEN_12275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12277 = 7'h4b == _myNewVec_33_T_3[6:0] ? myVec_75 : _GEN_12276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12278 = 7'h4c == _myNewVec_33_T_3[6:0] ? myVec_76 : _GEN_12277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12279 = 7'h4d == _myNewVec_33_T_3[6:0] ? myVec_77 : _GEN_12278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12280 = 7'h4e == _myNewVec_33_T_3[6:0] ? myVec_78 : _GEN_12279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12281 = 7'h4f == _myNewVec_33_T_3[6:0] ? myVec_79 : _GEN_12280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12282 = 7'h50 == _myNewVec_33_T_3[6:0] ? myVec_80 : _GEN_12281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12283 = 7'h51 == _myNewVec_33_T_3[6:0] ? myVec_81 : _GEN_12282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12284 = 7'h52 == _myNewVec_33_T_3[6:0] ? myVec_82 : _GEN_12283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12285 = 7'h53 == _myNewVec_33_T_3[6:0] ? myVec_83 : _GEN_12284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12286 = 7'h54 == _myNewVec_33_T_3[6:0] ? myVec_84 : _GEN_12285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12287 = 7'h55 == _myNewVec_33_T_3[6:0] ? myVec_85 : _GEN_12286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12288 = 7'h56 == _myNewVec_33_T_3[6:0] ? myVec_86 : _GEN_12287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12289 = 7'h57 == _myNewVec_33_T_3[6:0] ? myVec_87 : _GEN_12288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12290 = 7'h58 == _myNewVec_33_T_3[6:0] ? myVec_88 : _GEN_12289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12291 = 7'h59 == _myNewVec_33_T_3[6:0] ? myVec_89 : _GEN_12290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12292 = 7'h5a == _myNewVec_33_T_3[6:0] ? myVec_90 : _GEN_12291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12293 = 7'h5b == _myNewVec_33_T_3[6:0] ? myVec_91 : _GEN_12292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12294 = 7'h5c == _myNewVec_33_T_3[6:0] ? myVec_92 : _GEN_12293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12295 = 7'h5d == _myNewVec_33_T_3[6:0] ? myVec_93 : _GEN_12294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12296 = 7'h5e == _myNewVec_33_T_3[6:0] ? myVec_94 : _GEN_12295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12297 = 7'h5f == _myNewVec_33_T_3[6:0] ? myVec_95 : _GEN_12296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12298 = 7'h60 == _myNewVec_33_T_3[6:0] ? myVec_96 : _GEN_12297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12299 = 7'h61 == _myNewVec_33_T_3[6:0] ? myVec_97 : _GEN_12298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12300 = 7'h62 == _myNewVec_33_T_3[6:0] ? myVec_98 : _GEN_12299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12301 = 7'h63 == _myNewVec_33_T_3[6:0] ? myVec_99 : _GEN_12300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12302 = 7'h64 == _myNewVec_33_T_3[6:0] ? myVec_100 : _GEN_12301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12303 = 7'h65 == _myNewVec_33_T_3[6:0] ? myVec_101 : _GEN_12302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12304 = 7'h66 == _myNewVec_33_T_3[6:0] ? myVec_102 : _GEN_12303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12305 = 7'h67 == _myNewVec_33_T_3[6:0] ? myVec_103 : _GEN_12304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12306 = 7'h68 == _myNewVec_33_T_3[6:0] ? myVec_104 : _GEN_12305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12307 = 7'h69 == _myNewVec_33_T_3[6:0] ? myVec_105 : _GEN_12306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12308 = 7'h6a == _myNewVec_33_T_3[6:0] ? myVec_106 : _GEN_12307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12309 = 7'h6b == _myNewVec_33_T_3[6:0] ? myVec_107 : _GEN_12308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12310 = 7'h6c == _myNewVec_33_T_3[6:0] ? myVec_108 : _GEN_12309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12311 = 7'h6d == _myNewVec_33_T_3[6:0] ? myVec_109 : _GEN_12310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12312 = 7'h6e == _myNewVec_33_T_3[6:0] ? myVec_110 : _GEN_12311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12313 = 7'h6f == _myNewVec_33_T_3[6:0] ? myVec_111 : _GEN_12312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12314 = 7'h70 == _myNewVec_33_T_3[6:0] ? myVec_112 : _GEN_12313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12315 = 7'h71 == _myNewVec_33_T_3[6:0] ? myVec_113 : _GEN_12314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12316 = 7'h72 == _myNewVec_33_T_3[6:0] ? myVec_114 : _GEN_12315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12317 = 7'h73 == _myNewVec_33_T_3[6:0] ? myVec_115 : _GEN_12316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12318 = 7'h74 == _myNewVec_33_T_3[6:0] ? myVec_116 : _GEN_12317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12319 = 7'h75 == _myNewVec_33_T_3[6:0] ? myVec_117 : _GEN_12318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12320 = 7'h76 == _myNewVec_33_T_3[6:0] ? myVec_118 : _GEN_12319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12321 = 7'h77 == _myNewVec_33_T_3[6:0] ? myVec_119 : _GEN_12320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12322 = 7'h78 == _myNewVec_33_T_3[6:0] ? myVec_120 : _GEN_12321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12323 = 7'h79 == _myNewVec_33_T_3[6:0] ? myVec_121 : _GEN_12322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12324 = 7'h7a == _myNewVec_33_T_3[6:0] ? myVec_122 : _GEN_12323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12325 = 7'h7b == _myNewVec_33_T_3[6:0] ? myVec_123 : _GEN_12324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12326 = 7'h7c == _myNewVec_33_T_3[6:0] ? myVec_124 : _GEN_12325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12327 = 7'h7d == _myNewVec_33_T_3[6:0] ? myVec_125 : _GEN_12326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12328 = 7'h7e == _myNewVec_33_T_3[6:0] ? myVec_126 : _GEN_12327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_33 = 7'h7f == _myNewVec_33_T_3[6:0] ? myVec_127 : _GEN_12328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_32_T_3 = _myNewVec_127_T_1 + 16'h5f; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_12331 = 7'h1 == _myNewVec_32_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12332 = 7'h2 == _myNewVec_32_T_3[6:0] ? myVec_2 : _GEN_12331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12333 = 7'h3 == _myNewVec_32_T_3[6:0] ? myVec_3 : _GEN_12332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12334 = 7'h4 == _myNewVec_32_T_3[6:0] ? myVec_4 : _GEN_12333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12335 = 7'h5 == _myNewVec_32_T_3[6:0] ? myVec_5 : _GEN_12334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12336 = 7'h6 == _myNewVec_32_T_3[6:0] ? myVec_6 : _GEN_12335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12337 = 7'h7 == _myNewVec_32_T_3[6:0] ? myVec_7 : _GEN_12336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12338 = 7'h8 == _myNewVec_32_T_3[6:0] ? myVec_8 : _GEN_12337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12339 = 7'h9 == _myNewVec_32_T_3[6:0] ? myVec_9 : _GEN_12338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12340 = 7'ha == _myNewVec_32_T_3[6:0] ? myVec_10 : _GEN_12339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12341 = 7'hb == _myNewVec_32_T_3[6:0] ? myVec_11 : _GEN_12340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12342 = 7'hc == _myNewVec_32_T_3[6:0] ? myVec_12 : _GEN_12341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12343 = 7'hd == _myNewVec_32_T_3[6:0] ? myVec_13 : _GEN_12342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12344 = 7'he == _myNewVec_32_T_3[6:0] ? myVec_14 : _GEN_12343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12345 = 7'hf == _myNewVec_32_T_3[6:0] ? myVec_15 : _GEN_12344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12346 = 7'h10 == _myNewVec_32_T_3[6:0] ? myVec_16 : _GEN_12345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12347 = 7'h11 == _myNewVec_32_T_3[6:0] ? myVec_17 : _GEN_12346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12348 = 7'h12 == _myNewVec_32_T_3[6:0] ? myVec_18 : _GEN_12347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12349 = 7'h13 == _myNewVec_32_T_3[6:0] ? myVec_19 : _GEN_12348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12350 = 7'h14 == _myNewVec_32_T_3[6:0] ? myVec_20 : _GEN_12349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12351 = 7'h15 == _myNewVec_32_T_3[6:0] ? myVec_21 : _GEN_12350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12352 = 7'h16 == _myNewVec_32_T_3[6:0] ? myVec_22 : _GEN_12351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12353 = 7'h17 == _myNewVec_32_T_3[6:0] ? myVec_23 : _GEN_12352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12354 = 7'h18 == _myNewVec_32_T_3[6:0] ? myVec_24 : _GEN_12353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12355 = 7'h19 == _myNewVec_32_T_3[6:0] ? myVec_25 : _GEN_12354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12356 = 7'h1a == _myNewVec_32_T_3[6:0] ? myVec_26 : _GEN_12355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12357 = 7'h1b == _myNewVec_32_T_3[6:0] ? myVec_27 : _GEN_12356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12358 = 7'h1c == _myNewVec_32_T_3[6:0] ? myVec_28 : _GEN_12357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12359 = 7'h1d == _myNewVec_32_T_3[6:0] ? myVec_29 : _GEN_12358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12360 = 7'h1e == _myNewVec_32_T_3[6:0] ? myVec_30 : _GEN_12359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12361 = 7'h1f == _myNewVec_32_T_3[6:0] ? myVec_31 : _GEN_12360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12362 = 7'h20 == _myNewVec_32_T_3[6:0] ? myVec_32 : _GEN_12361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12363 = 7'h21 == _myNewVec_32_T_3[6:0] ? myVec_33 : _GEN_12362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12364 = 7'h22 == _myNewVec_32_T_3[6:0] ? myVec_34 : _GEN_12363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12365 = 7'h23 == _myNewVec_32_T_3[6:0] ? myVec_35 : _GEN_12364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12366 = 7'h24 == _myNewVec_32_T_3[6:0] ? myVec_36 : _GEN_12365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12367 = 7'h25 == _myNewVec_32_T_3[6:0] ? myVec_37 : _GEN_12366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12368 = 7'h26 == _myNewVec_32_T_3[6:0] ? myVec_38 : _GEN_12367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12369 = 7'h27 == _myNewVec_32_T_3[6:0] ? myVec_39 : _GEN_12368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12370 = 7'h28 == _myNewVec_32_T_3[6:0] ? myVec_40 : _GEN_12369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12371 = 7'h29 == _myNewVec_32_T_3[6:0] ? myVec_41 : _GEN_12370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12372 = 7'h2a == _myNewVec_32_T_3[6:0] ? myVec_42 : _GEN_12371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12373 = 7'h2b == _myNewVec_32_T_3[6:0] ? myVec_43 : _GEN_12372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12374 = 7'h2c == _myNewVec_32_T_3[6:0] ? myVec_44 : _GEN_12373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12375 = 7'h2d == _myNewVec_32_T_3[6:0] ? myVec_45 : _GEN_12374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12376 = 7'h2e == _myNewVec_32_T_3[6:0] ? myVec_46 : _GEN_12375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12377 = 7'h2f == _myNewVec_32_T_3[6:0] ? myVec_47 : _GEN_12376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12378 = 7'h30 == _myNewVec_32_T_3[6:0] ? myVec_48 : _GEN_12377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12379 = 7'h31 == _myNewVec_32_T_3[6:0] ? myVec_49 : _GEN_12378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12380 = 7'h32 == _myNewVec_32_T_3[6:0] ? myVec_50 : _GEN_12379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12381 = 7'h33 == _myNewVec_32_T_3[6:0] ? myVec_51 : _GEN_12380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12382 = 7'h34 == _myNewVec_32_T_3[6:0] ? myVec_52 : _GEN_12381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12383 = 7'h35 == _myNewVec_32_T_3[6:0] ? myVec_53 : _GEN_12382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12384 = 7'h36 == _myNewVec_32_T_3[6:0] ? myVec_54 : _GEN_12383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12385 = 7'h37 == _myNewVec_32_T_3[6:0] ? myVec_55 : _GEN_12384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12386 = 7'h38 == _myNewVec_32_T_3[6:0] ? myVec_56 : _GEN_12385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12387 = 7'h39 == _myNewVec_32_T_3[6:0] ? myVec_57 : _GEN_12386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12388 = 7'h3a == _myNewVec_32_T_3[6:0] ? myVec_58 : _GEN_12387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12389 = 7'h3b == _myNewVec_32_T_3[6:0] ? myVec_59 : _GEN_12388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12390 = 7'h3c == _myNewVec_32_T_3[6:0] ? myVec_60 : _GEN_12389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12391 = 7'h3d == _myNewVec_32_T_3[6:0] ? myVec_61 : _GEN_12390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12392 = 7'h3e == _myNewVec_32_T_3[6:0] ? myVec_62 : _GEN_12391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12393 = 7'h3f == _myNewVec_32_T_3[6:0] ? myVec_63 : _GEN_12392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12394 = 7'h40 == _myNewVec_32_T_3[6:0] ? myVec_64 : _GEN_12393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12395 = 7'h41 == _myNewVec_32_T_3[6:0] ? myVec_65 : _GEN_12394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12396 = 7'h42 == _myNewVec_32_T_3[6:0] ? myVec_66 : _GEN_12395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12397 = 7'h43 == _myNewVec_32_T_3[6:0] ? myVec_67 : _GEN_12396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12398 = 7'h44 == _myNewVec_32_T_3[6:0] ? myVec_68 : _GEN_12397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12399 = 7'h45 == _myNewVec_32_T_3[6:0] ? myVec_69 : _GEN_12398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12400 = 7'h46 == _myNewVec_32_T_3[6:0] ? myVec_70 : _GEN_12399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12401 = 7'h47 == _myNewVec_32_T_3[6:0] ? myVec_71 : _GEN_12400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12402 = 7'h48 == _myNewVec_32_T_3[6:0] ? myVec_72 : _GEN_12401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12403 = 7'h49 == _myNewVec_32_T_3[6:0] ? myVec_73 : _GEN_12402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12404 = 7'h4a == _myNewVec_32_T_3[6:0] ? myVec_74 : _GEN_12403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12405 = 7'h4b == _myNewVec_32_T_3[6:0] ? myVec_75 : _GEN_12404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12406 = 7'h4c == _myNewVec_32_T_3[6:0] ? myVec_76 : _GEN_12405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12407 = 7'h4d == _myNewVec_32_T_3[6:0] ? myVec_77 : _GEN_12406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12408 = 7'h4e == _myNewVec_32_T_3[6:0] ? myVec_78 : _GEN_12407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12409 = 7'h4f == _myNewVec_32_T_3[6:0] ? myVec_79 : _GEN_12408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12410 = 7'h50 == _myNewVec_32_T_3[6:0] ? myVec_80 : _GEN_12409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12411 = 7'h51 == _myNewVec_32_T_3[6:0] ? myVec_81 : _GEN_12410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12412 = 7'h52 == _myNewVec_32_T_3[6:0] ? myVec_82 : _GEN_12411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12413 = 7'h53 == _myNewVec_32_T_3[6:0] ? myVec_83 : _GEN_12412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12414 = 7'h54 == _myNewVec_32_T_3[6:0] ? myVec_84 : _GEN_12413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12415 = 7'h55 == _myNewVec_32_T_3[6:0] ? myVec_85 : _GEN_12414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12416 = 7'h56 == _myNewVec_32_T_3[6:0] ? myVec_86 : _GEN_12415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12417 = 7'h57 == _myNewVec_32_T_3[6:0] ? myVec_87 : _GEN_12416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12418 = 7'h58 == _myNewVec_32_T_3[6:0] ? myVec_88 : _GEN_12417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12419 = 7'h59 == _myNewVec_32_T_3[6:0] ? myVec_89 : _GEN_12418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12420 = 7'h5a == _myNewVec_32_T_3[6:0] ? myVec_90 : _GEN_12419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12421 = 7'h5b == _myNewVec_32_T_3[6:0] ? myVec_91 : _GEN_12420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12422 = 7'h5c == _myNewVec_32_T_3[6:0] ? myVec_92 : _GEN_12421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12423 = 7'h5d == _myNewVec_32_T_3[6:0] ? myVec_93 : _GEN_12422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12424 = 7'h5e == _myNewVec_32_T_3[6:0] ? myVec_94 : _GEN_12423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12425 = 7'h5f == _myNewVec_32_T_3[6:0] ? myVec_95 : _GEN_12424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12426 = 7'h60 == _myNewVec_32_T_3[6:0] ? myVec_96 : _GEN_12425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12427 = 7'h61 == _myNewVec_32_T_3[6:0] ? myVec_97 : _GEN_12426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12428 = 7'h62 == _myNewVec_32_T_3[6:0] ? myVec_98 : _GEN_12427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12429 = 7'h63 == _myNewVec_32_T_3[6:0] ? myVec_99 : _GEN_12428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12430 = 7'h64 == _myNewVec_32_T_3[6:0] ? myVec_100 : _GEN_12429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12431 = 7'h65 == _myNewVec_32_T_3[6:0] ? myVec_101 : _GEN_12430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12432 = 7'h66 == _myNewVec_32_T_3[6:0] ? myVec_102 : _GEN_12431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12433 = 7'h67 == _myNewVec_32_T_3[6:0] ? myVec_103 : _GEN_12432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12434 = 7'h68 == _myNewVec_32_T_3[6:0] ? myVec_104 : _GEN_12433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12435 = 7'h69 == _myNewVec_32_T_3[6:0] ? myVec_105 : _GEN_12434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12436 = 7'h6a == _myNewVec_32_T_3[6:0] ? myVec_106 : _GEN_12435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12437 = 7'h6b == _myNewVec_32_T_3[6:0] ? myVec_107 : _GEN_12436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12438 = 7'h6c == _myNewVec_32_T_3[6:0] ? myVec_108 : _GEN_12437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12439 = 7'h6d == _myNewVec_32_T_3[6:0] ? myVec_109 : _GEN_12438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12440 = 7'h6e == _myNewVec_32_T_3[6:0] ? myVec_110 : _GEN_12439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12441 = 7'h6f == _myNewVec_32_T_3[6:0] ? myVec_111 : _GEN_12440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12442 = 7'h70 == _myNewVec_32_T_3[6:0] ? myVec_112 : _GEN_12441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12443 = 7'h71 == _myNewVec_32_T_3[6:0] ? myVec_113 : _GEN_12442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12444 = 7'h72 == _myNewVec_32_T_3[6:0] ? myVec_114 : _GEN_12443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12445 = 7'h73 == _myNewVec_32_T_3[6:0] ? myVec_115 : _GEN_12444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12446 = 7'h74 == _myNewVec_32_T_3[6:0] ? myVec_116 : _GEN_12445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12447 = 7'h75 == _myNewVec_32_T_3[6:0] ? myVec_117 : _GEN_12446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12448 = 7'h76 == _myNewVec_32_T_3[6:0] ? myVec_118 : _GEN_12447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12449 = 7'h77 == _myNewVec_32_T_3[6:0] ? myVec_119 : _GEN_12448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12450 = 7'h78 == _myNewVec_32_T_3[6:0] ? myVec_120 : _GEN_12449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12451 = 7'h79 == _myNewVec_32_T_3[6:0] ? myVec_121 : _GEN_12450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12452 = 7'h7a == _myNewVec_32_T_3[6:0] ? myVec_122 : _GEN_12451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12453 = 7'h7b == _myNewVec_32_T_3[6:0] ? myVec_123 : _GEN_12452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12454 = 7'h7c == _myNewVec_32_T_3[6:0] ? myVec_124 : _GEN_12453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12455 = 7'h7d == _myNewVec_32_T_3[6:0] ? myVec_125 : _GEN_12454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12456 = 7'h7e == _myNewVec_32_T_3[6:0] ? myVec_126 : _GEN_12455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_32 = 7'h7f == _myNewVec_32_T_3[6:0] ? myVec_127 : _GEN_12456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [255:0] myNewWire_lo_hi_lo_lo = {myNewVec_39,myNewVec_38,myNewVec_37,myNewVec_36,myNewVec_35,myNewVec_34,
    myNewVec_33,myNewVec_32}; // @[hh_datapath_chisel.scala 238:27]
  wire [511:0] myNewWire_lo_hi_lo = {myNewVec_47,myNewVec_46,myNewVec_45,myNewVec_44,myNewVec_43,myNewVec_42,myNewVec_41
    ,myNewVec_40,myNewWire_lo_hi_lo_lo}; // @[hh_datapath_chisel.scala 238:27]
  wire [1023:0] myNewWire_lo_hi = {myNewVec_63,myNewVec_62,myNewVec_61,myNewVec_60,myNewVec_59,myNewVec_58,myNewVec_57,
    myNewVec_56,myNewWire_lo_hi_hi_lo,myNewWire_lo_hi_lo}; // @[hh_datapath_chisel.scala 238:27]
  wire [15:0] _myNewVec_31_T_3 = _myNewVec_127_T_1 + 16'h60; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_12459 = 7'h1 == _myNewVec_31_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12460 = 7'h2 == _myNewVec_31_T_3[6:0] ? myVec_2 : _GEN_12459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12461 = 7'h3 == _myNewVec_31_T_3[6:0] ? myVec_3 : _GEN_12460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12462 = 7'h4 == _myNewVec_31_T_3[6:0] ? myVec_4 : _GEN_12461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12463 = 7'h5 == _myNewVec_31_T_3[6:0] ? myVec_5 : _GEN_12462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12464 = 7'h6 == _myNewVec_31_T_3[6:0] ? myVec_6 : _GEN_12463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12465 = 7'h7 == _myNewVec_31_T_3[6:0] ? myVec_7 : _GEN_12464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12466 = 7'h8 == _myNewVec_31_T_3[6:0] ? myVec_8 : _GEN_12465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12467 = 7'h9 == _myNewVec_31_T_3[6:0] ? myVec_9 : _GEN_12466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12468 = 7'ha == _myNewVec_31_T_3[6:0] ? myVec_10 : _GEN_12467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12469 = 7'hb == _myNewVec_31_T_3[6:0] ? myVec_11 : _GEN_12468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12470 = 7'hc == _myNewVec_31_T_3[6:0] ? myVec_12 : _GEN_12469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12471 = 7'hd == _myNewVec_31_T_3[6:0] ? myVec_13 : _GEN_12470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12472 = 7'he == _myNewVec_31_T_3[6:0] ? myVec_14 : _GEN_12471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12473 = 7'hf == _myNewVec_31_T_3[6:0] ? myVec_15 : _GEN_12472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12474 = 7'h10 == _myNewVec_31_T_3[6:0] ? myVec_16 : _GEN_12473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12475 = 7'h11 == _myNewVec_31_T_3[6:0] ? myVec_17 : _GEN_12474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12476 = 7'h12 == _myNewVec_31_T_3[6:0] ? myVec_18 : _GEN_12475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12477 = 7'h13 == _myNewVec_31_T_3[6:0] ? myVec_19 : _GEN_12476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12478 = 7'h14 == _myNewVec_31_T_3[6:0] ? myVec_20 : _GEN_12477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12479 = 7'h15 == _myNewVec_31_T_3[6:0] ? myVec_21 : _GEN_12478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12480 = 7'h16 == _myNewVec_31_T_3[6:0] ? myVec_22 : _GEN_12479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12481 = 7'h17 == _myNewVec_31_T_3[6:0] ? myVec_23 : _GEN_12480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12482 = 7'h18 == _myNewVec_31_T_3[6:0] ? myVec_24 : _GEN_12481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12483 = 7'h19 == _myNewVec_31_T_3[6:0] ? myVec_25 : _GEN_12482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12484 = 7'h1a == _myNewVec_31_T_3[6:0] ? myVec_26 : _GEN_12483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12485 = 7'h1b == _myNewVec_31_T_3[6:0] ? myVec_27 : _GEN_12484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12486 = 7'h1c == _myNewVec_31_T_3[6:0] ? myVec_28 : _GEN_12485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12487 = 7'h1d == _myNewVec_31_T_3[6:0] ? myVec_29 : _GEN_12486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12488 = 7'h1e == _myNewVec_31_T_3[6:0] ? myVec_30 : _GEN_12487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12489 = 7'h1f == _myNewVec_31_T_3[6:0] ? myVec_31 : _GEN_12488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12490 = 7'h20 == _myNewVec_31_T_3[6:0] ? myVec_32 : _GEN_12489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12491 = 7'h21 == _myNewVec_31_T_3[6:0] ? myVec_33 : _GEN_12490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12492 = 7'h22 == _myNewVec_31_T_3[6:0] ? myVec_34 : _GEN_12491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12493 = 7'h23 == _myNewVec_31_T_3[6:0] ? myVec_35 : _GEN_12492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12494 = 7'h24 == _myNewVec_31_T_3[6:0] ? myVec_36 : _GEN_12493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12495 = 7'h25 == _myNewVec_31_T_3[6:0] ? myVec_37 : _GEN_12494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12496 = 7'h26 == _myNewVec_31_T_3[6:0] ? myVec_38 : _GEN_12495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12497 = 7'h27 == _myNewVec_31_T_3[6:0] ? myVec_39 : _GEN_12496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12498 = 7'h28 == _myNewVec_31_T_3[6:0] ? myVec_40 : _GEN_12497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12499 = 7'h29 == _myNewVec_31_T_3[6:0] ? myVec_41 : _GEN_12498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12500 = 7'h2a == _myNewVec_31_T_3[6:0] ? myVec_42 : _GEN_12499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12501 = 7'h2b == _myNewVec_31_T_3[6:0] ? myVec_43 : _GEN_12500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12502 = 7'h2c == _myNewVec_31_T_3[6:0] ? myVec_44 : _GEN_12501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12503 = 7'h2d == _myNewVec_31_T_3[6:0] ? myVec_45 : _GEN_12502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12504 = 7'h2e == _myNewVec_31_T_3[6:0] ? myVec_46 : _GEN_12503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12505 = 7'h2f == _myNewVec_31_T_3[6:0] ? myVec_47 : _GEN_12504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12506 = 7'h30 == _myNewVec_31_T_3[6:0] ? myVec_48 : _GEN_12505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12507 = 7'h31 == _myNewVec_31_T_3[6:0] ? myVec_49 : _GEN_12506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12508 = 7'h32 == _myNewVec_31_T_3[6:0] ? myVec_50 : _GEN_12507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12509 = 7'h33 == _myNewVec_31_T_3[6:0] ? myVec_51 : _GEN_12508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12510 = 7'h34 == _myNewVec_31_T_3[6:0] ? myVec_52 : _GEN_12509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12511 = 7'h35 == _myNewVec_31_T_3[6:0] ? myVec_53 : _GEN_12510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12512 = 7'h36 == _myNewVec_31_T_3[6:0] ? myVec_54 : _GEN_12511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12513 = 7'h37 == _myNewVec_31_T_3[6:0] ? myVec_55 : _GEN_12512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12514 = 7'h38 == _myNewVec_31_T_3[6:0] ? myVec_56 : _GEN_12513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12515 = 7'h39 == _myNewVec_31_T_3[6:0] ? myVec_57 : _GEN_12514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12516 = 7'h3a == _myNewVec_31_T_3[6:0] ? myVec_58 : _GEN_12515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12517 = 7'h3b == _myNewVec_31_T_3[6:0] ? myVec_59 : _GEN_12516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12518 = 7'h3c == _myNewVec_31_T_3[6:0] ? myVec_60 : _GEN_12517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12519 = 7'h3d == _myNewVec_31_T_3[6:0] ? myVec_61 : _GEN_12518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12520 = 7'h3e == _myNewVec_31_T_3[6:0] ? myVec_62 : _GEN_12519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12521 = 7'h3f == _myNewVec_31_T_3[6:0] ? myVec_63 : _GEN_12520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12522 = 7'h40 == _myNewVec_31_T_3[6:0] ? myVec_64 : _GEN_12521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12523 = 7'h41 == _myNewVec_31_T_3[6:0] ? myVec_65 : _GEN_12522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12524 = 7'h42 == _myNewVec_31_T_3[6:0] ? myVec_66 : _GEN_12523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12525 = 7'h43 == _myNewVec_31_T_3[6:0] ? myVec_67 : _GEN_12524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12526 = 7'h44 == _myNewVec_31_T_3[6:0] ? myVec_68 : _GEN_12525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12527 = 7'h45 == _myNewVec_31_T_3[6:0] ? myVec_69 : _GEN_12526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12528 = 7'h46 == _myNewVec_31_T_3[6:0] ? myVec_70 : _GEN_12527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12529 = 7'h47 == _myNewVec_31_T_3[6:0] ? myVec_71 : _GEN_12528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12530 = 7'h48 == _myNewVec_31_T_3[6:0] ? myVec_72 : _GEN_12529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12531 = 7'h49 == _myNewVec_31_T_3[6:0] ? myVec_73 : _GEN_12530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12532 = 7'h4a == _myNewVec_31_T_3[6:0] ? myVec_74 : _GEN_12531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12533 = 7'h4b == _myNewVec_31_T_3[6:0] ? myVec_75 : _GEN_12532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12534 = 7'h4c == _myNewVec_31_T_3[6:0] ? myVec_76 : _GEN_12533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12535 = 7'h4d == _myNewVec_31_T_3[6:0] ? myVec_77 : _GEN_12534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12536 = 7'h4e == _myNewVec_31_T_3[6:0] ? myVec_78 : _GEN_12535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12537 = 7'h4f == _myNewVec_31_T_3[6:0] ? myVec_79 : _GEN_12536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12538 = 7'h50 == _myNewVec_31_T_3[6:0] ? myVec_80 : _GEN_12537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12539 = 7'h51 == _myNewVec_31_T_3[6:0] ? myVec_81 : _GEN_12538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12540 = 7'h52 == _myNewVec_31_T_3[6:0] ? myVec_82 : _GEN_12539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12541 = 7'h53 == _myNewVec_31_T_3[6:0] ? myVec_83 : _GEN_12540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12542 = 7'h54 == _myNewVec_31_T_3[6:0] ? myVec_84 : _GEN_12541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12543 = 7'h55 == _myNewVec_31_T_3[6:0] ? myVec_85 : _GEN_12542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12544 = 7'h56 == _myNewVec_31_T_3[6:0] ? myVec_86 : _GEN_12543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12545 = 7'h57 == _myNewVec_31_T_3[6:0] ? myVec_87 : _GEN_12544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12546 = 7'h58 == _myNewVec_31_T_3[6:0] ? myVec_88 : _GEN_12545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12547 = 7'h59 == _myNewVec_31_T_3[6:0] ? myVec_89 : _GEN_12546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12548 = 7'h5a == _myNewVec_31_T_3[6:0] ? myVec_90 : _GEN_12547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12549 = 7'h5b == _myNewVec_31_T_3[6:0] ? myVec_91 : _GEN_12548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12550 = 7'h5c == _myNewVec_31_T_3[6:0] ? myVec_92 : _GEN_12549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12551 = 7'h5d == _myNewVec_31_T_3[6:0] ? myVec_93 : _GEN_12550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12552 = 7'h5e == _myNewVec_31_T_3[6:0] ? myVec_94 : _GEN_12551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12553 = 7'h5f == _myNewVec_31_T_3[6:0] ? myVec_95 : _GEN_12552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12554 = 7'h60 == _myNewVec_31_T_3[6:0] ? myVec_96 : _GEN_12553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12555 = 7'h61 == _myNewVec_31_T_3[6:0] ? myVec_97 : _GEN_12554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12556 = 7'h62 == _myNewVec_31_T_3[6:0] ? myVec_98 : _GEN_12555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12557 = 7'h63 == _myNewVec_31_T_3[6:0] ? myVec_99 : _GEN_12556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12558 = 7'h64 == _myNewVec_31_T_3[6:0] ? myVec_100 : _GEN_12557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12559 = 7'h65 == _myNewVec_31_T_3[6:0] ? myVec_101 : _GEN_12558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12560 = 7'h66 == _myNewVec_31_T_3[6:0] ? myVec_102 : _GEN_12559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12561 = 7'h67 == _myNewVec_31_T_3[6:0] ? myVec_103 : _GEN_12560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12562 = 7'h68 == _myNewVec_31_T_3[6:0] ? myVec_104 : _GEN_12561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12563 = 7'h69 == _myNewVec_31_T_3[6:0] ? myVec_105 : _GEN_12562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12564 = 7'h6a == _myNewVec_31_T_3[6:0] ? myVec_106 : _GEN_12563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12565 = 7'h6b == _myNewVec_31_T_3[6:0] ? myVec_107 : _GEN_12564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12566 = 7'h6c == _myNewVec_31_T_3[6:0] ? myVec_108 : _GEN_12565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12567 = 7'h6d == _myNewVec_31_T_3[6:0] ? myVec_109 : _GEN_12566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12568 = 7'h6e == _myNewVec_31_T_3[6:0] ? myVec_110 : _GEN_12567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12569 = 7'h6f == _myNewVec_31_T_3[6:0] ? myVec_111 : _GEN_12568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12570 = 7'h70 == _myNewVec_31_T_3[6:0] ? myVec_112 : _GEN_12569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12571 = 7'h71 == _myNewVec_31_T_3[6:0] ? myVec_113 : _GEN_12570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12572 = 7'h72 == _myNewVec_31_T_3[6:0] ? myVec_114 : _GEN_12571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12573 = 7'h73 == _myNewVec_31_T_3[6:0] ? myVec_115 : _GEN_12572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12574 = 7'h74 == _myNewVec_31_T_3[6:0] ? myVec_116 : _GEN_12573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12575 = 7'h75 == _myNewVec_31_T_3[6:0] ? myVec_117 : _GEN_12574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12576 = 7'h76 == _myNewVec_31_T_3[6:0] ? myVec_118 : _GEN_12575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12577 = 7'h77 == _myNewVec_31_T_3[6:0] ? myVec_119 : _GEN_12576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12578 = 7'h78 == _myNewVec_31_T_3[6:0] ? myVec_120 : _GEN_12577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12579 = 7'h79 == _myNewVec_31_T_3[6:0] ? myVec_121 : _GEN_12578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12580 = 7'h7a == _myNewVec_31_T_3[6:0] ? myVec_122 : _GEN_12579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12581 = 7'h7b == _myNewVec_31_T_3[6:0] ? myVec_123 : _GEN_12580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12582 = 7'h7c == _myNewVec_31_T_3[6:0] ? myVec_124 : _GEN_12581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12583 = 7'h7d == _myNewVec_31_T_3[6:0] ? myVec_125 : _GEN_12582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12584 = 7'h7e == _myNewVec_31_T_3[6:0] ? myVec_126 : _GEN_12583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_31 = 7'h7f == _myNewVec_31_T_3[6:0] ? myVec_127 : _GEN_12584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_30_T_3 = _myNewVec_127_T_1 + 16'h61; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_12587 = 7'h1 == _myNewVec_30_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12588 = 7'h2 == _myNewVec_30_T_3[6:0] ? myVec_2 : _GEN_12587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12589 = 7'h3 == _myNewVec_30_T_3[6:0] ? myVec_3 : _GEN_12588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12590 = 7'h4 == _myNewVec_30_T_3[6:0] ? myVec_4 : _GEN_12589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12591 = 7'h5 == _myNewVec_30_T_3[6:0] ? myVec_5 : _GEN_12590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12592 = 7'h6 == _myNewVec_30_T_3[6:0] ? myVec_6 : _GEN_12591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12593 = 7'h7 == _myNewVec_30_T_3[6:0] ? myVec_7 : _GEN_12592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12594 = 7'h8 == _myNewVec_30_T_3[6:0] ? myVec_8 : _GEN_12593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12595 = 7'h9 == _myNewVec_30_T_3[6:0] ? myVec_9 : _GEN_12594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12596 = 7'ha == _myNewVec_30_T_3[6:0] ? myVec_10 : _GEN_12595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12597 = 7'hb == _myNewVec_30_T_3[6:0] ? myVec_11 : _GEN_12596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12598 = 7'hc == _myNewVec_30_T_3[6:0] ? myVec_12 : _GEN_12597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12599 = 7'hd == _myNewVec_30_T_3[6:0] ? myVec_13 : _GEN_12598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12600 = 7'he == _myNewVec_30_T_3[6:0] ? myVec_14 : _GEN_12599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12601 = 7'hf == _myNewVec_30_T_3[6:0] ? myVec_15 : _GEN_12600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12602 = 7'h10 == _myNewVec_30_T_3[6:0] ? myVec_16 : _GEN_12601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12603 = 7'h11 == _myNewVec_30_T_3[6:0] ? myVec_17 : _GEN_12602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12604 = 7'h12 == _myNewVec_30_T_3[6:0] ? myVec_18 : _GEN_12603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12605 = 7'h13 == _myNewVec_30_T_3[6:0] ? myVec_19 : _GEN_12604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12606 = 7'h14 == _myNewVec_30_T_3[6:0] ? myVec_20 : _GEN_12605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12607 = 7'h15 == _myNewVec_30_T_3[6:0] ? myVec_21 : _GEN_12606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12608 = 7'h16 == _myNewVec_30_T_3[6:0] ? myVec_22 : _GEN_12607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12609 = 7'h17 == _myNewVec_30_T_3[6:0] ? myVec_23 : _GEN_12608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12610 = 7'h18 == _myNewVec_30_T_3[6:0] ? myVec_24 : _GEN_12609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12611 = 7'h19 == _myNewVec_30_T_3[6:0] ? myVec_25 : _GEN_12610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12612 = 7'h1a == _myNewVec_30_T_3[6:0] ? myVec_26 : _GEN_12611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12613 = 7'h1b == _myNewVec_30_T_3[6:0] ? myVec_27 : _GEN_12612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12614 = 7'h1c == _myNewVec_30_T_3[6:0] ? myVec_28 : _GEN_12613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12615 = 7'h1d == _myNewVec_30_T_3[6:0] ? myVec_29 : _GEN_12614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12616 = 7'h1e == _myNewVec_30_T_3[6:0] ? myVec_30 : _GEN_12615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12617 = 7'h1f == _myNewVec_30_T_3[6:0] ? myVec_31 : _GEN_12616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12618 = 7'h20 == _myNewVec_30_T_3[6:0] ? myVec_32 : _GEN_12617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12619 = 7'h21 == _myNewVec_30_T_3[6:0] ? myVec_33 : _GEN_12618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12620 = 7'h22 == _myNewVec_30_T_3[6:0] ? myVec_34 : _GEN_12619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12621 = 7'h23 == _myNewVec_30_T_3[6:0] ? myVec_35 : _GEN_12620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12622 = 7'h24 == _myNewVec_30_T_3[6:0] ? myVec_36 : _GEN_12621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12623 = 7'h25 == _myNewVec_30_T_3[6:0] ? myVec_37 : _GEN_12622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12624 = 7'h26 == _myNewVec_30_T_3[6:0] ? myVec_38 : _GEN_12623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12625 = 7'h27 == _myNewVec_30_T_3[6:0] ? myVec_39 : _GEN_12624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12626 = 7'h28 == _myNewVec_30_T_3[6:0] ? myVec_40 : _GEN_12625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12627 = 7'h29 == _myNewVec_30_T_3[6:0] ? myVec_41 : _GEN_12626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12628 = 7'h2a == _myNewVec_30_T_3[6:0] ? myVec_42 : _GEN_12627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12629 = 7'h2b == _myNewVec_30_T_3[6:0] ? myVec_43 : _GEN_12628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12630 = 7'h2c == _myNewVec_30_T_3[6:0] ? myVec_44 : _GEN_12629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12631 = 7'h2d == _myNewVec_30_T_3[6:0] ? myVec_45 : _GEN_12630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12632 = 7'h2e == _myNewVec_30_T_3[6:0] ? myVec_46 : _GEN_12631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12633 = 7'h2f == _myNewVec_30_T_3[6:0] ? myVec_47 : _GEN_12632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12634 = 7'h30 == _myNewVec_30_T_3[6:0] ? myVec_48 : _GEN_12633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12635 = 7'h31 == _myNewVec_30_T_3[6:0] ? myVec_49 : _GEN_12634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12636 = 7'h32 == _myNewVec_30_T_3[6:0] ? myVec_50 : _GEN_12635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12637 = 7'h33 == _myNewVec_30_T_3[6:0] ? myVec_51 : _GEN_12636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12638 = 7'h34 == _myNewVec_30_T_3[6:0] ? myVec_52 : _GEN_12637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12639 = 7'h35 == _myNewVec_30_T_3[6:0] ? myVec_53 : _GEN_12638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12640 = 7'h36 == _myNewVec_30_T_3[6:0] ? myVec_54 : _GEN_12639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12641 = 7'h37 == _myNewVec_30_T_3[6:0] ? myVec_55 : _GEN_12640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12642 = 7'h38 == _myNewVec_30_T_3[6:0] ? myVec_56 : _GEN_12641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12643 = 7'h39 == _myNewVec_30_T_3[6:0] ? myVec_57 : _GEN_12642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12644 = 7'h3a == _myNewVec_30_T_3[6:0] ? myVec_58 : _GEN_12643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12645 = 7'h3b == _myNewVec_30_T_3[6:0] ? myVec_59 : _GEN_12644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12646 = 7'h3c == _myNewVec_30_T_3[6:0] ? myVec_60 : _GEN_12645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12647 = 7'h3d == _myNewVec_30_T_3[6:0] ? myVec_61 : _GEN_12646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12648 = 7'h3e == _myNewVec_30_T_3[6:0] ? myVec_62 : _GEN_12647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12649 = 7'h3f == _myNewVec_30_T_3[6:0] ? myVec_63 : _GEN_12648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12650 = 7'h40 == _myNewVec_30_T_3[6:0] ? myVec_64 : _GEN_12649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12651 = 7'h41 == _myNewVec_30_T_3[6:0] ? myVec_65 : _GEN_12650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12652 = 7'h42 == _myNewVec_30_T_3[6:0] ? myVec_66 : _GEN_12651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12653 = 7'h43 == _myNewVec_30_T_3[6:0] ? myVec_67 : _GEN_12652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12654 = 7'h44 == _myNewVec_30_T_3[6:0] ? myVec_68 : _GEN_12653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12655 = 7'h45 == _myNewVec_30_T_3[6:0] ? myVec_69 : _GEN_12654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12656 = 7'h46 == _myNewVec_30_T_3[6:0] ? myVec_70 : _GEN_12655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12657 = 7'h47 == _myNewVec_30_T_3[6:0] ? myVec_71 : _GEN_12656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12658 = 7'h48 == _myNewVec_30_T_3[6:0] ? myVec_72 : _GEN_12657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12659 = 7'h49 == _myNewVec_30_T_3[6:0] ? myVec_73 : _GEN_12658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12660 = 7'h4a == _myNewVec_30_T_3[6:0] ? myVec_74 : _GEN_12659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12661 = 7'h4b == _myNewVec_30_T_3[6:0] ? myVec_75 : _GEN_12660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12662 = 7'h4c == _myNewVec_30_T_3[6:0] ? myVec_76 : _GEN_12661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12663 = 7'h4d == _myNewVec_30_T_3[6:0] ? myVec_77 : _GEN_12662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12664 = 7'h4e == _myNewVec_30_T_3[6:0] ? myVec_78 : _GEN_12663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12665 = 7'h4f == _myNewVec_30_T_3[6:0] ? myVec_79 : _GEN_12664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12666 = 7'h50 == _myNewVec_30_T_3[6:0] ? myVec_80 : _GEN_12665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12667 = 7'h51 == _myNewVec_30_T_3[6:0] ? myVec_81 : _GEN_12666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12668 = 7'h52 == _myNewVec_30_T_3[6:0] ? myVec_82 : _GEN_12667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12669 = 7'h53 == _myNewVec_30_T_3[6:0] ? myVec_83 : _GEN_12668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12670 = 7'h54 == _myNewVec_30_T_3[6:0] ? myVec_84 : _GEN_12669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12671 = 7'h55 == _myNewVec_30_T_3[6:0] ? myVec_85 : _GEN_12670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12672 = 7'h56 == _myNewVec_30_T_3[6:0] ? myVec_86 : _GEN_12671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12673 = 7'h57 == _myNewVec_30_T_3[6:0] ? myVec_87 : _GEN_12672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12674 = 7'h58 == _myNewVec_30_T_3[6:0] ? myVec_88 : _GEN_12673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12675 = 7'h59 == _myNewVec_30_T_3[6:0] ? myVec_89 : _GEN_12674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12676 = 7'h5a == _myNewVec_30_T_3[6:0] ? myVec_90 : _GEN_12675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12677 = 7'h5b == _myNewVec_30_T_3[6:0] ? myVec_91 : _GEN_12676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12678 = 7'h5c == _myNewVec_30_T_3[6:0] ? myVec_92 : _GEN_12677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12679 = 7'h5d == _myNewVec_30_T_3[6:0] ? myVec_93 : _GEN_12678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12680 = 7'h5e == _myNewVec_30_T_3[6:0] ? myVec_94 : _GEN_12679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12681 = 7'h5f == _myNewVec_30_T_3[6:0] ? myVec_95 : _GEN_12680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12682 = 7'h60 == _myNewVec_30_T_3[6:0] ? myVec_96 : _GEN_12681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12683 = 7'h61 == _myNewVec_30_T_3[6:0] ? myVec_97 : _GEN_12682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12684 = 7'h62 == _myNewVec_30_T_3[6:0] ? myVec_98 : _GEN_12683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12685 = 7'h63 == _myNewVec_30_T_3[6:0] ? myVec_99 : _GEN_12684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12686 = 7'h64 == _myNewVec_30_T_3[6:0] ? myVec_100 : _GEN_12685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12687 = 7'h65 == _myNewVec_30_T_3[6:0] ? myVec_101 : _GEN_12686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12688 = 7'h66 == _myNewVec_30_T_3[6:0] ? myVec_102 : _GEN_12687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12689 = 7'h67 == _myNewVec_30_T_3[6:0] ? myVec_103 : _GEN_12688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12690 = 7'h68 == _myNewVec_30_T_3[6:0] ? myVec_104 : _GEN_12689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12691 = 7'h69 == _myNewVec_30_T_3[6:0] ? myVec_105 : _GEN_12690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12692 = 7'h6a == _myNewVec_30_T_3[6:0] ? myVec_106 : _GEN_12691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12693 = 7'h6b == _myNewVec_30_T_3[6:0] ? myVec_107 : _GEN_12692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12694 = 7'h6c == _myNewVec_30_T_3[6:0] ? myVec_108 : _GEN_12693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12695 = 7'h6d == _myNewVec_30_T_3[6:0] ? myVec_109 : _GEN_12694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12696 = 7'h6e == _myNewVec_30_T_3[6:0] ? myVec_110 : _GEN_12695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12697 = 7'h6f == _myNewVec_30_T_3[6:0] ? myVec_111 : _GEN_12696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12698 = 7'h70 == _myNewVec_30_T_3[6:0] ? myVec_112 : _GEN_12697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12699 = 7'h71 == _myNewVec_30_T_3[6:0] ? myVec_113 : _GEN_12698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12700 = 7'h72 == _myNewVec_30_T_3[6:0] ? myVec_114 : _GEN_12699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12701 = 7'h73 == _myNewVec_30_T_3[6:0] ? myVec_115 : _GEN_12700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12702 = 7'h74 == _myNewVec_30_T_3[6:0] ? myVec_116 : _GEN_12701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12703 = 7'h75 == _myNewVec_30_T_3[6:0] ? myVec_117 : _GEN_12702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12704 = 7'h76 == _myNewVec_30_T_3[6:0] ? myVec_118 : _GEN_12703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12705 = 7'h77 == _myNewVec_30_T_3[6:0] ? myVec_119 : _GEN_12704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12706 = 7'h78 == _myNewVec_30_T_3[6:0] ? myVec_120 : _GEN_12705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12707 = 7'h79 == _myNewVec_30_T_3[6:0] ? myVec_121 : _GEN_12706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12708 = 7'h7a == _myNewVec_30_T_3[6:0] ? myVec_122 : _GEN_12707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12709 = 7'h7b == _myNewVec_30_T_3[6:0] ? myVec_123 : _GEN_12708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12710 = 7'h7c == _myNewVec_30_T_3[6:0] ? myVec_124 : _GEN_12709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12711 = 7'h7d == _myNewVec_30_T_3[6:0] ? myVec_125 : _GEN_12710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12712 = 7'h7e == _myNewVec_30_T_3[6:0] ? myVec_126 : _GEN_12711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_30 = 7'h7f == _myNewVec_30_T_3[6:0] ? myVec_127 : _GEN_12712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_29_T_3 = _myNewVec_127_T_1 + 16'h62; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_12715 = 7'h1 == _myNewVec_29_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12716 = 7'h2 == _myNewVec_29_T_3[6:0] ? myVec_2 : _GEN_12715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12717 = 7'h3 == _myNewVec_29_T_3[6:0] ? myVec_3 : _GEN_12716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12718 = 7'h4 == _myNewVec_29_T_3[6:0] ? myVec_4 : _GEN_12717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12719 = 7'h5 == _myNewVec_29_T_3[6:0] ? myVec_5 : _GEN_12718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12720 = 7'h6 == _myNewVec_29_T_3[6:0] ? myVec_6 : _GEN_12719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12721 = 7'h7 == _myNewVec_29_T_3[6:0] ? myVec_7 : _GEN_12720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12722 = 7'h8 == _myNewVec_29_T_3[6:0] ? myVec_8 : _GEN_12721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12723 = 7'h9 == _myNewVec_29_T_3[6:0] ? myVec_9 : _GEN_12722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12724 = 7'ha == _myNewVec_29_T_3[6:0] ? myVec_10 : _GEN_12723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12725 = 7'hb == _myNewVec_29_T_3[6:0] ? myVec_11 : _GEN_12724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12726 = 7'hc == _myNewVec_29_T_3[6:0] ? myVec_12 : _GEN_12725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12727 = 7'hd == _myNewVec_29_T_3[6:0] ? myVec_13 : _GEN_12726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12728 = 7'he == _myNewVec_29_T_3[6:0] ? myVec_14 : _GEN_12727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12729 = 7'hf == _myNewVec_29_T_3[6:0] ? myVec_15 : _GEN_12728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12730 = 7'h10 == _myNewVec_29_T_3[6:0] ? myVec_16 : _GEN_12729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12731 = 7'h11 == _myNewVec_29_T_3[6:0] ? myVec_17 : _GEN_12730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12732 = 7'h12 == _myNewVec_29_T_3[6:0] ? myVec_18 : _GEN_12731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12733 = 7'h13 == _myNewVec_29_T_3[6:0] ? myVec_19 : _GEN_12732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12734 = 7'h14 == _myNewVec_29_T_3[6:0] ? myVec_20 : _GEN_12733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12735 = 7'h15 == _myNewVec_29_T_3[6:0] ? myVec_21 : _GEN_12734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12736 = 7'h16 == _myNewVec_29_T_3[6:0] ? myVec_22 : _GEN_12735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12737 = 7'h17 == _myNewVec_29_T_3[6:0] ? myVec_23 : _GEN_12736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12738 = 7'h18 == _myNewVec_29_T_3[6:0] ? myVec_24 : _GEN_12737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12739 = 7'h19 == _myNewVec_29_T_3[6:0] ? myVec_25 : _GEN_12738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12740 = 7'h1a == _myNewVec_29_T_3[6:0] ? myVec_26 : _GEN_12739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12741 = 7'h1b == _myNewVec_29_T_3[6:0] ? myVec_27 : _GEN_12740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12742 = 7'h1c == _myNewVec_29_T_3[6:0] ? myVec_28 : _GEN_12741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12743 = 7'h1d == _myNewVec_29_T_3[6:0] ? myVec_29 : _GEN_12742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12744 = 7'h1e == _myNewVec_29_T_3[6:0] ? myVec_30 : _GEN_12743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12745 = 7'h1f == _myNewVec_29_T_3[6:0] ? myVec_31 : _GEN_12744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12746 = 7'h20 == _myNewVec_29_T_3[6:0] ? myVec_32 : _GEN_12745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12747 = 7'h21 == _myNewVec_29_T_3[6:0] ? myVec_33 : _GEN_12746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12748 = 7'h22 == _myNewVec_29_T_3[6:0] ? myVec_34 : _GEN_12747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12749 = 7'h23 == _myNewVec_29_T_3[6:0] ? myVec_35 : _GEN_12748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12750 = 7'h24 == _myNewVec_29_T_3[6:0] ? myVec_36 : _GEN_12749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12751 = 7'h25 == _myNewVec_29_T_3[6:0] ? myVec_37 : _GEN_12750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12752 = 7'h26 == _myNewVec_29_T_3[6:0] ? myVec_38 : _GEN_12751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12753 = 7'h27 == _myNewVec_29_T_3[6:0] ? myVec_39 : _GEN_12752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12754 = 7'h28 == _myNewVec_29_T_3[6:0] ? myVec_40 : _GEN_12753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12755 = 7'h29 == _myNewVec_29_T_3[6:0] ? myVec_41 : _GEN_12754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12756 = 7'h2a == _myNewVec_29_T_3[6:0] ? myVec_42 : _GEN_12755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12757 = 7'h2b == _myNewVec_29_T_3[6:0] ? myVec_43 : _GEN_12756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12758 = 7'h2c == _myNewVec_29_T_3[6:0] ? myVec_44 : _GEN_12757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12759 = 7'h2d == _myNewVec_29_T_3[6:0] ? myVec_45 : _GEN_12758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12760 = 7'h2e == _myNewVec_29_T_3[6:0] ? myVec_46 : _GEN_12759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12761 = 7'h2f == _myNewVec_29_T_3[6:0] ? myVec_47 : _GEN_12760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12762 = 7'h30 == _myNewVec_29_T_3[6:0] ? myVec_48 : _GEN_12761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12763 = 7'h31 == _myNewVec_29_T_3[6:0] ? myVec_49 : _GEN_12762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12764 = 7'h32 == _myNewVec_29_T_3[6:0] ? myVec_50 : _GEN_12763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12765 = 7'h33 == _myNewVec_29_T_3[6:0] ? myVec_51 : _GEN_12764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12766 = 7'h34 == _myNewVec_29_T_3[6:0] ? myVec_52 : _GEN_12765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12767 = 7'h35 == _myNewVec_29_T_3[6:0] ? myVec_53 : _GEN_12766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12768 = 7'h36 == _myNewVec_29_T_3[6:0] ? myVec_54 : _GEN_12767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12769 = 7'h37 == _myNewVec_29_T_3[6:0] ? myVec_55 : _GEN_12768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12770 = 7'h38 == _myNewVec_29_T_3[6:0] ? myVec_56 : _GEN_12769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12771 = 7'h39 == _myNewVec_29_T_3[6:0] ? myVec_57 : _GEN_12770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12772 = 7'h3a == _myNewVec_29_T_3[6:0] ? myVec_58 : _GEN_12771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12773 = 7'h3b == _myNewVec_29_T_3[6:0] ? myVec_59 : _GEN_12772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12774 = 7'h3c == _myNewVec_29_T_3[6:0] ? myVec_60 : _GEN_12773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12775 = 7'h3d == _myNewVec_29_T_3[6:0] ? myVec_61 : _GEN_12774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12776 = 7'h3e == _myNewVec_29_T_3[6:0] ? myVec_62 : _GEN_12775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12777 = 7'h3f == _myNewVec_29_T_3[6:0] ? myVec_63 : _GEN_12776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12778 = 7'h40 == _myNewVec_29_T_3[6:0] ? myVec_64 : _GEN_12777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12779 = 7'h41 == _myNewVec_29_T_3[6:0] ? myVec_65 : _GEN_12778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12780 = 7'h42 == _myNewVec_29_T_3[6:0] ? myVec_66 : _GEN_12779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12781 = 7'h43 == _myNewVec_29_T_3[6:0] ? myVec_67 : _GEN_12780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12782 = 7'h44 == _myNewVec_29_T_3[6:0] ? myVec_68 : _GEN_12781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12783 = 7'h45 == _myNewVec_29_T_3[6:0] ? myVec_69 : _GEN_12782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12784 = 7'h46 == _myNewVec_29_T_3[6:0] ? myVec_70 : _GEN_12783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12785 = 7'h47 == _myNewVec_29_T_3[6:0] ? myVec_71 : _GEN_12784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12786 = 7'h48 == _myNewVec_29_T_3[6:0] ? myVec_72 : _GEN_12785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12787 = 7'h49 == _myNewVec_29_T_3[6:0] ? myVec_73 : _GEN_12786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12788 = 7'h4a == _myNewVec_29_T_3[6:0] ? myVec_74 : _GEN_12787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12789 = 7'h4b == _myNewVec_29_T_3[6:0] ? myVec_75 : _GEN_12788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12790 = 7'h4c == _myNewVec_29_T_3[6:0] ? myVec_76 : _GEN_12789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12791 = 7'h4d == _myNewVec_29_T_3[6:0] ? myVec_77 : _GEN_12790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12792 = 7'h4e == _myNewVec_29_T_3[6:0] ? myVec_78 : _GEN_12791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12793 = 7'h4f == _myNewVec_29_T_3[6:0] ? myVec_79 : _GEN_12792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12794 = 7'h50 == _myNewVec_29_T_3[6:0] ? myVec_80 : _GEN_12793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12795 = 7'h51 == _myNewVec_29_T_3[6:0] ? myVec_81 : _GEN_12794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12796 = 7'h52 == _myNewVec_29_T_3[6:0] ? myVec_82 : _GEN_12795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12797 = 7'h53 == _myNewVec_29_T_3[6:0] ? myVec_83 : _GEN_12796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12798 = 7'h54 == _myNewVec_29_T_3[6:0] ? myVec_84 : _GEN_12797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12799 = 7'h55 == _myNewVec_29_T_3[6:0] ? myVec_85 : _GEN_12798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12800 = 7'h56 == _myNewVec_29_T_3[6:0] ? myVec_86 : _GEN_12799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12801 = 7'h57 == _myNewVec_29_T_3[6:0] ? myVec_87 : _GEN_12800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12802 = 7'h58 == _myNewVec_29_T_3[6:0] ? myVec_88 : _GEN_12801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12803 = 7'h59 == _myNewVec_29_T_3[6:0] ? myVec_89 : _GEN_12802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12804 = 7'h5a == _myNewVec_29_T_3[6:0] ? myVec_90 : _GEN_12803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12805 = 7'h5b == _myNewVec_29_T_3[6:0] ? myVec_91 : _GEN_12804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12806 = 7'h5c == _myNewVec_29_T_3[6:0] ? myVec_92 : _GEN_12805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12807 = 7'h5d == _myNewVec_29_T_3[6:0] ? myVec_93 : _GEN_12806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12808 = 7'h5e == _myNewVec_29_T_3[6:0] ? myVec_94 : _GEN_12807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12809 = 7'h5f == _myNewVec_29_T_3[6:0] ? myVec_95 : _GEN_12808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12810 = 7'h60 == _myNewVec_29_T_3[6:0] ? myVec_96 : _GEN_12809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12811 = 7'h61 == _myNewVec_29_T_3[6:0] ? myVec_97 : _GEN_12810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12812 = 7'h62 == _myNewVec_29_T_3[6:0] ? myVec_98 : _GEN_12811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12813 = 7'h63 == _myNewVec_29_T_3[6:0] ? myVec_99 : _GEN_12812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12814 = 7'h64 == _myNewVec_29_T_3[6:0] ? myVec_100 : _GEN_12813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12815 = 7'h65 == _myNewVec_29_T_3[6:0] ? myVec_101 : _GEN_12814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12816 = 7'h66 == _myNewVec_29_T_3[6:0] ? myVec_102 : _GEN_12815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12817 = 7'h67 == _myNewVec_29_T_3[6:0] ? myVec_103 : _GEN_12816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12818 = 7'h68 == _myNewVec_29_T_3[6:0] ? myVec_104 : _GEN_12817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12819 = 7'h69 == _myNewVec_29_T_3[6:0] ? myVec_105 : _GEN_12818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12820 = 7'h6a == _myNewVec_29_T_3[6:0] ? myVec_106 : _GEN_12819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12821 = 7'h6b == _myNewVec_29_T_3[6:0] ? myVec_107 : _GEN_12820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12822 = 7'h6c == _myNewVec_29_T_3[6:0] ? myVec_108 : _GEN_12821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12823 = 7'h6d == _myNewVec_29_T_3[6:0] ? myVec_109 : _GEN_12822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12824 = 7'h6e == _myNewVec_29_T_3[6:0] ? myVec_110 : _GEN_12823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12825 = 7'h6f == _myNewVec_29_T_3[6:0] ? myVec_111 : _GEN_12824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12826 = 7'h70 == _myNewVec_29_T_3[6:0] ? myVec_112 : _GEN_12825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12827 = 7'h71 == _myNewVec_29_T_3[6:0] ? myVec_113 : _GEN_12826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12828 = 7'h72 == _myNewVec_29_T_3[6:0] ? myVec_114 : _GEN_12827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12829 = 7'h73 == _myNewVec_29_T_3[6:0] ? myVec_115 : _GEN_12828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12830 = 7'h74 == _myNewVec_29_T_3[6:0] ? myVec_116 : _GEN_12829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12831 = 7'h75 == _myNewVec_29_T_3[6:0] ? myVec_117 : _GEN_12830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12832 = 7'h76 == _myNewVec_29_T_3[6:0] ? myVec_118 : _GEN_12831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12833 = 7'h77 == _myNewVec_29_T_3[6:0] ? myVec_119 : _GEN_12832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12834 = 7'h78 == _myNewVec_29_T_3[6:0] ? myVec_120 : _GEN_12833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12835 = 7'h79 == _myNewVec_29_T_3[6:0] ? myVec_121 : _GEN_12834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12836 = 7'h7a == _myNewVec_29_T_3[6:0] ? myVec_122 : _GEN_12835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12837 = 7'h7b == _myNewVec_29_T_3[6:0] ? myVec_123 : _GEN_12836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12838 = 7'h7c == _myNewVec_29_T_3[6:0] ? myVec_124 : _GEN_12837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12839 = 7'h7d == _myNewVec_29_T_3[6:0] ? myVec_125 : _GEN_12838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12840 = 7'h7e == _myNewVec_29_T_3[6:0] ? myVec_126 : _GEN_12839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_29 = 7'h7f == _myNewVec_29_T_3[6:0] ? myVec_127 : _GEN_12840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_28_T_3 = _myNewVec_127_T_1 + 16'h63; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_12843 = 7'h1 == _myNewVec_28_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12844 = 7'h2 == _myNewVec_28_T_3[6:0] ? myVec_2 : _GEN_12843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12845 = 7'h3 == _myNewVec_28_T_3[6:0] ? myVec_3 : _GEN_12844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12846 = 7'h4 == _myNewVec_28_T_3[6:0] ? myVec_4 : _GEN_12845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12847 = 7'h5 == _myNewVec_28_T_3[6:0] ? myVec_5 : _GEN_12846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12848 = 7'h6 == _myNewVec_28_T_3[6:0] ? myVec_6 : _GEN_12847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12849 = 7'h7 == _myNewVec_28_T_3[6:0] ? myVec_7 : _GEN_12848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12850 = 7'h8 == _myNewVec_28_T_3[6:0] ? myVec_8 : _GEN_12849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12851 = 7'h9 == _myNewVec_28_T_3[6:0] ? myVec_9 : _GEN_12850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12852 = 7'ha == _myNewVec_28_T_3[6:0] ? myVec_10 : _GEN_12851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12853 = 7'hb == _myNewVec_28_T_3[6:0] ? myVec_11 : _GEN_12852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12854 = 7'hc == _myNewVec_28_T_3[6:0] ? myVec_12 : _GEN_12853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12855 = 7'hd == _myNewVec_28_T_3[6:0] ? myVec_13 : _GEN_12854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12856 = 7'he == _myNewVec_28_T_3[6:0] ? myVec_14 : _GEN_12855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12857 = 7'hf == _myNewVec_28_T_3[6:0] ? myVec_15 : _GEN_12856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12858 = 7'h10 == _myNewVec_28_T_3[6:0] ? myVec_16 : _GEN_12857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12859 = 7'h11 == _myNewVec_28_T_3[6:0] ? myVec_17 : _GEN_12858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12860 = 7'h12 == _myNewVec_28_T_3[6:0] ? myVec_18 : _GEN_12859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12861 = 7'h13 == _myNewVec_28_T_3[6:0] ? myVec_19 : _GEN_12860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12862 = 7'h14 == _myNewVec_28_T_3[6:0] ? myVec_20 : _GEN_12861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12863 = 7'h15 == _myNewVec_28_T_3[6:0] ? myVec_21 : _GEN_12862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12864 = 7'h16 == _myNewVec_28_T_3[6:0] ? myVec_22 : _GEN_12863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12865 = 7'h17 == _myNewVec_28_T_3[6:0] ? myVec_23 : _GEN_12864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12866 = 7'h18 == _myNewVec_28_T_3[6:0] ? myVec_24 : _GEN_12865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12867 = 7'h19 == _myNewVec_28_T_3[6:0] ? myVec_25 : _GEN_12866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12868 = 7'h1a == _myNewVec_28_T_3[6:0] ? myVec_26 : _GEN_12867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12869 = 7'h1b == _myNewVec_28_T_3[6:0] ? myVec_27 : _GEN_12868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12870 = 7'h1c == _myNewVec_28_T_3[6:0] ? myVec_28 : _GEN_12869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12871 = 7'h1d == _myNewVec_28_T_3[6:0] ? myVec_29 : _GEN_12870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12872 = 7'h1e == _myNewVec_28_T_3[6:0] ? myVec_30 : _GEN_12871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12873 = 7'h1f == _myNewVec_28_T_3[6:0] ? myVec_31 : _GEN_12872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12874 = 7'h20 == _myNewVec_28_T_3[6:0] ? myVec_32 : _GEN_12873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12875 = 7'h21 == _myNewVec_28_T_3[6:0] ? myVec_33 : _GEN_12874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12876 = 7'h22 == _myNewVec_28_T_3[6:0] ? myVec_34 : _GEN_12875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12877 = 7'h23 == _myNewVec_28_T_3[6:0] ? myVec_35 : _GEN_12876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12878 = 7'h24 == _myNewVec_28_T_3[6:0] ? myVec_36 : _GEN_12877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12879 = 7'h25 == _myNewVec_28_T_3[6:0] ? myVec_37 : _GEN_12878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12880 = 7'h26 == _myNewVec_28_T_3[6:0] ? myVec_38 : _GEN_12879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12881 = 7'h27 == _myNewVec_28_T_3[6:0] ? myVec_39 : _GEN_12880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12882 = 7'h28 == _myNewVec_28_T_3[6:0] ? myVec_40 : _GEN_12881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12883 = 7'h29 == _myNewVec_28_T_3[6:0] ? myVec_41 : _GEN_12882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12884 = 7'h2a == _myNewVec_28_T_3[6:0] ? myVec_42 : _GEN_12883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12885 = 7'h2b == _myNewVec_28_T_3[6:0] ? myVec_43 : _GEN_12884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12886 = 7'h2c == _myNewVec_28_T_3[6:0] ? myVec_44 : _GEN_12885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12887 = 7'h2d == _myNewVec_28_T_3[6:0] ? myVec_45 : _GEN_12886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12888 = 7'h2e == _myNewVec_28_T_3[6:0] ? myVec_46 : _GEN_12887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12889 = 7'h2f == _myNewVec_28_T_3[6:0] ? myVec_47 : _GEN_12888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12890 = 7'h30 == _myNewVec_28_T_3[6:0] ? myVec_48 : _GEN_12889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12891 = 7'h31 == _myNewVec_28_T_3[6:0] ? myVec_49 : _GEN_12890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12892 = 7'h32 == _myNewVec_28_T_3[6:0] ? myVec_50 : _GEN_12891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12893 = 7'h33 == _myNewVec_28_T_3[6:0] ? myVec_51 : _GEN_12892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12894 = 7'h34 == _myNewVec_28_T_3[6:0] ? myVec_52 : _GEN_12893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12895 = 7'h35 == _myNewVec_28_T_3[6:0] ? myVec_53 : _GEN_12894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12896 = 7'h36 == _myNewVec_28_T_3[6:0] ? myVec_54 : _GEN_12895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12897 = 7'h37 == _myNewVec_28_T_3[6:0] ? myVec_55 : _GEN_12896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12898 = 7'h38 == _myNewVec_28_T_3[6:0] ? myVec_56 : _GEN_12897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12899 = 7'h39 == _myNewVec_28_T_3[6:0] ? myVec_57 : _GEN_12898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12900 = 7'h3a == _myNewVec_28_T_3[6:0] ? myVec_58 : _GEN_12899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12901 = 7'h3b == _myNewVec_28_T_3[6:0] ? myVec_59 : _GEN_12900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12902 = 7'h3c == _myNewVec_28_T_3[6:0] ? myVec_60 : _GEN_12901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12903 = 7'h3d == _myNewVec_28_T_3[6:0] ? myVec_61 : _GEN_12902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12904 = 7'h3e == _myNewVec_28_T_3[6:0] ? myVec_62 : _GEN_12903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12905 = 7'h3f == _myNewVec_28_T_3[6:0] ? myVec_63 : _GEN_12904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12906 = 7'h40 == _myNewVec_28_T_3[6:0] ? myVec_64 : _GEN_12905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12907 = 7'h41 == _myNewVec_28_T_3[6:0] ? myVec_65 : _GEN_12906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12908 = 7'h42 == _myNewVec_28_T_3[6:0] ? myVec_66 : _GEN_12907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12909 = 7'h43 == _myNewVec_28_T_3[6:0] ? myVec_67 : _GEN_12908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12910 = 7'h44 == _myNewVec_28_T_3[6:0] ? myVec_68 : _GEN_12909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12911 = 7'h45 == _myNewVec_28_T_3[6:0] ? myVec_69 : _GEN_12910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12912 = 7'h46 == _myNewVec_28_T_3[6:0] ? myVec_70 : _GEN_12911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12913 = 7'h47 == _myNewVec_28_T_3[6:0] ? myVec_71 : _GEN_12912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12914 = 7'h48 == _myNewVec_28_T_3[6:0] ? myVec_72 : _GEN_12913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12915 = 7'h49 == _myNewVec_28_T_3[6:0] ? myVec_73 : _GEN_12914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12916 = 7'h4a == _myNewVec_28_T_3[6:0] ? myVec_74 : _GEN_12915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12917 = 7'h4b == _myNewVec_28_T_3[6:0] ? myVec_75 : _GEN_12916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12918 = 7'h4c == _myNewVec_28_T_3[6:0] ? myVec_76 : _GEN_12917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12919 = 7'h4d == _myNewVec_28_T_3[6:0] ? myVec_77 : _GEN_12918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12920 = 7'h4e == _myNewVec_28_T_3[6:0] ? myVec_78 : _GEN_12919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12921 = 7'h4f == _myNewVec_28_T_3[6:0] ? myVec_79 : _GEN_12920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12922 = 7'h50 == _myNewVec_28_T_3[6:0] ? myVec_80 : _GEN_12921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12923 = 7'h51 == _myNewVec_28_T_3[6:0] ? myVec_81 : _GEN_12922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12924 = 7'h52 == _myNewVec_28_T_3[6:0] ? myVec_82 : _GEN_12923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12925 = 7'h53 == _myNewVec_28_T_3[6:0] ? myVec_83 : _GEN_12924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12926 = 7'h54 == _myNewVec_28_T_3[6:0] ? myVec_84 : _GEN_12925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12927 = 7'h55 == _myNewVec_28_T_3[6:0] ? myVec_85 : _GEN_12926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12928 = 7'h56 == _myNewVec_28_T_3[6:0] ? myVec_86 : _GEN_12927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12929 = 7'h57 == _myNewVec_28_T_3[6:0] ? myVec_87 : _GEN_12928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12930 = 7'h58 == _myNewVec_28_T_3[6:0] ? myVec_88 : _GEN_12929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12931 = 7'h59 == _myNewVec_28_T_3[6:0] ? myVec_89 : _GEN_12930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12932 = 7'h5a == _myNewVec_28_T_3[6:0] ? myVec_90 : _GEN_12931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12933 = 7'h5b == _myNewVec_28_T_3[6:0] ? myVec_91 : _GEN_12932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12934 = 7'h5c == _myNewVec_28_T_3[6:0] ? myVec_92 : _GEN_12933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12935 = 7'h5d == _myNewVec_28_T_3[6:0] ? myVec_93 : _GEN_12934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12936 = 7'h5e == _myNewVec_28_T_3[6:0] ? myVec_94 : _GEN_12935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12937 = 7'h5f == _myNewVec_28_T_3[6:0] ? myVec_95 : _GEN_12936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12938 = 7'h60 == _myNewVec_28_T_3[6:0] ? myVec_96 : _GEN_12937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12939 = 7'h61 == _myNewVec_28_T_3[6:0] ? myVec_97 : _GEN_12938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12940 = 7'h62 == _myNewVec_28_T_3[6:0] ? myVec_98 : _GEN_12939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12941 = 7'h63 == _myNewVec_28_T_3[6:0] ? myVec_99 : _GEN_12940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12942 = 7'h64 == _myNewVec_28_T_3[6:0] ? myVec_100 : _GEN_12941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12943 = 7'h65 == _myNewVec_28_T_3[6:0] ? myVec_101 : _GEN_12942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12944 = 7'h66 == _myNewVec_28_T_3[6:0] ? myVec_102 : _GEN_12943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12945 = 7'h67 == _myNewVec_28_T_3[6:0] ? myVec_103 : _GEN_12944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12946 = 7'h68 == _myNewVec_28_T_3[6:0] ? myVec_104 : _GEN_12945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12947 = 7'h69 == _myNewVec_28_T_3[6:0] ? myVec_105 : _GEN_12946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12948 = 7'h6a == _myNewVec_28_T_3[6:0] ? myVec_106 : _GEN_12947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12949 = 7'h6b == _myNewVec_28_T_3[6:0] ? myVec_107 : _GEN_12948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12950 = 7'h6c == _myNewVec_28_T_3[6:0] ? myVec_108 : _GEN_12949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12951 = 7'h6d == _myNewVec_28_T_3[6:0] ? myVec_109 : _GEN_12950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12952 = 7'h6e == _myNewVec_28_T_3[6:0] ? myVec_110 : _GEN_12951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12953 = 7'h6f == _myNewVec_28_T_3[6:0] ? myVec_111 : _GEN_12952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12954 = 7'h70 == _myNewVec_28_T_3[6:0] ? myVec_112 : _GEN_12953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12955 = 7'h71 == _myNewVec_28_T_3[6:0] ? myVec_113 : _GEN_12954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12956 = 7'h72 == _myNewVec_28_T_3[6:0] ? myVec_114 : _GEN_12955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12957 = 7'h73 == _myNewVec_28_T_3[6:0] ? myVec_115 : _GEN_12956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12958 = 7'h74 == _myNewVec_28_T_3[6:0] ? myVec_116 : _GEN_12957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12959 = 7'h75 == _myNewVec_28_T_3[6:0] ? myVec_117 : _GEN_12958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12960 = 7'h76 == _myNewVec_28_T_3[6:0] ? myVec_118 : _GEN_12959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12961 = 7'h77 == _myNewVec_28_T_3[6:0] ? myVec_119 : _GEN_12960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12962 = 7'h78 == _myNewVec_28_T_3[6:0] ? myVec_120 : _GEN_12961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12963 = 7'h79 == _myNewVec_28_T_3[6:0] ? myVec_121 : _GEN_12962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12964 = 7'h7a == _myNewVec_28_T_3[6:0] ? myVec_122 : _GEN_12963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12965 = 7'h7b == _myNewVec_28_T_3[6:0] ? myVec_123 : _GEN_12964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12966 = 7'h7c == _myNewVec_28_T_3[6:0] ? myVec_124 : _GEN_12965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12967 = 7'h7d == _myNewVec_28_T_3[6:0] ? myVec_125 : _GEN_12966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12968 = 7'h7e == _myNewVec_28_T_3[6:0] ? myVec_126 : _GEN_12967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_28 = 7'h7f == _myNewVec_28_T_3[6:0] ? myVec_127 : _GEN_12968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_27_T_3 = _myNewVec_127_T_1 + 16'h64; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_12971 = 7'h1 == _myNewVec_27_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12972 = 7'h2 == _myNewVec_27_T_3[6:0] ? myVec_2 : _GEN_12971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12973 = 7'h3 == _myNewVec_27_T_3[6:0] ? myVec_3 : _GEN_12972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12974 = 7'h4 == _myNewVec_27_T_3[6:0] ? myVec_4 : _GEN_12973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12975 = 7'h5 == _myNewVec_27_T_3[6:0] ? myVec_5 : _GEN_12974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12976 = 7'h6 == _myNewVec_27_T_3[6:0] ? myVec_6 : _GEN_12975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12977 = 7'h7 == _myNewVec_27_T_3[6:0] ? myVec_7 : _GEN_12976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12978 = 7'h8 == _myNewVec_27_T_3[6:0] ? myVec_8 : _GEN_12977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12979 = 7'h9 == _myNewVec_27_T_3[6:0] ? myVec_9 : _GEN_12978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12980 = 7'ha == _myNewVec_27_T_3[6:0] ? myVec_10 : _GEN_12979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12981 = 7'hb == _myNewVec_27_T_3[6:0] ? myVec_11 : _GEN_12980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12982 = 7'hc == _myNewVec_27_T_3[6:0] ? myVec_12 : _GEN_12981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12983 = 7'hd == _myNewVec_27_T_3[6:0] ? myVec_13 : _GEN_12982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12984 = 7'he == _myNewVec_27_T_3[6:0] ? myVec_14 : _GEN_12983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12985 = 7'hf == _myNewVec_27_T_3[6:0] ? myVec_15 : _GEN_12984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12986 = 7'h10 == _myNewVec_27_T_3[6:0] ? myVec_16 : _GEN_12985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12987 = 7'h11 == _myNewVec_27_T_3[6:0] ? myVec_17 : _GEN_12986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12988 = 7'h12 == _myNewVec_27_T_3[6:0] ? myVec_18 : _GEN_12987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12989 = 7'h13 == _myNewVec_27_T_3[6:0] ? myVec_19 : _GEN_12988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12990 = 7'h14 == _myNewVec_27_T_3[6:0] ? myVec_20 : _GEN_12989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12991 = 7'h15 == _myNewVec_27_T_3[6:0] ? myVec_21 : _GEN_12990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12992 = 7'h16 == _myNewVec_27_T_3[6:0] ? myVec_22 : _GEN_12991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12993 = 7'h17 == _myNewVec_27_T_3[6:0] ? myVec_23 : _GEN_12992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12994 = 7'h18 == _myNewVec_27_T_3[6:0] ? myVec_24 : _GEN_12993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12995 = 7'h19 == _myNewVec_27_T_3[6:0] ? myVec_25 : _GEN_12994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12996 = 7'h1a == _myNewVec_27_T_3[6:0] ? myVec_26 : _GEN_12995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12997 = 7'h1b == _myNewVec_27_T_3[6:0] ? myVec_27 : _GEN_12996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12998 = 7'h1c == _myNewVec_27_T_3[6:0] ? myVec_28 : _GEN_12997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_12999 = 7'h1d == _myNewVec_27_T_3[6:0] ? myVec_29 : _GEN_12998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13000 = 7'h1e == _myNewVec_27_T_3[6:0] ? myVec_30 : _GEN_12999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13001 = 7'h1f == _myNewVec_27_T_3[6:0] ? myVec_31 : _GEN_13000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13002 = 7'h20 == _myNewVec_27_T_3[6:0] ? myVec_32 : _GEN_13001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13003 = 7'h21 == _myNewVec_27_T_3[6:0] ? myVec_33 : _GEN_13002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13004 = 7'h22 == _myNewVec_27_T_3[6:0] ? myVec_34 : _GEN_13003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13005 = 7'h23 == _myNewVec_27_T_3[6:0] ? myVec_35 : _GEN_13004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13006 = 7'h24 == _myNewVec_27_T_3[6:0] ? myVec_36 : _GEN_13005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13007 = 7'h25 == _myNewVec_27_T_3[6:0] ? myVec_37 : _GEN_13006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13008 = 7'h26 == _myNewVec_27_T_3[6:0] ? myVec_38 : _GEN_13007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13009 = 7'h27 == _myNewVec_27_T_3[6:0] ? myVec_39 : _GEN_13008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13010 = 7'h28 == _myNewVec_27_T_3[6:0] ? myVec_40 : _GEN_13009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13011 = 7'h29 == _myNewVec_27_T_3[6:0] ? myVec_41 : _GEN_13010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13012 = 7'h2a == _myNewVec_27_T_3[6:0] ? myVec_42 : _GEN_13011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13013 = 7'h2b == _myNewVec_27_T_3[6:0] ? myVec_43 : _GEN_13012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13014 = 7'h2c == _myNewVec_27_T_3[6:0] ? myVec_44 : _GEN_13013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13015 = 7'h2d == _myNewVec_27_T_3[6:0] ? myVec_45 : _GEN_13014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13016 = 7'h2e == _myNewVec_27_T_3[6:0] ? myVec_46 : _GEN_13015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13017 = 7'h2f == _myNewVec_27_T_3[6:0] ? myVec_47 : _GEN_13016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13018 = 7'h30 == _myNewVec_27_T_3[6:0] ? myVec_48 : _GEN_13017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13019 = 7'h31 == _myNewVec_27_T_3[6:0] ? myVec_49 : _GEN_13018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13020 = 7'h32 == _myNewVec_27_T_3[6:0] ? myVec_50 : _GEN_13019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13021 = 7'h33 == _myNewVec_27_T_3[6:0] ? myVec_51 : _GEN_13020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13022 = 7'h34 == _myNewVec_27_T_3[6:0] ? myVec_52 : _GEN_13021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13023 = 7'h35 == _myNewVec_27_T_3[6:0] ? myVec_53 : _GEN_13022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13024 = 7'h36 == _myNewVec_27_T_3[6:0] ? myVec_54 : _GEN_13023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13025 = 7'h37 == _myNewVec_27_T_3[6:0] ? myVec_55 : _GEN_13024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13026 = 7'h38 == _myNewVec_27_T_3[6:0] ? myVec_56 : _GEN_13025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13027 = 7'h39 == _myNewVec_27_T_3[6:0] ? myVec_57 : _GEN_13026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13028 = 7'h3a == _myNewVec_27_T_3[6:0] ? myVec_58 : _GEN_13027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13029 = 7'h3b == _myNewVec_27_T_3[6:0] ? myVec_59 : _GEN_13028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13030 = 7'h3c == _myNewVec_27_T_3[6:0] ? myVec_60 : _GEN_13029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13031 = 7'h3d == _myNewVec_27_T_3[6:0] ? myVec_61 : _GEN_13030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13032 = 7'h3e == _myNewVec_27_T_3[6:0] ? myVec_62 : _GEN_13031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13033 = 7'h3f == _myNewVec_27_T_3[6:0] ? myVec_63 : _GEN_13032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13034 = 7'h40 == _myNewVec_27_T_3[6:0] ? myVec_64 : _GEN_13033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13035 = 7'h41 == _myNewVec_27_T_3[6:0] ? myVec_65 : _GEN_13034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13036 = 7'h42 == _myNewVec_27_T_3[6:0] ? myVec_66 : _GEN_13035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13037 = 7'h43 == _myNewVec_27_T_3[6:0] ? myVec_67 : _GEN_13036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13038 = 7'h44 == _myNewVec_27_T_3[6:0] ? myVec_68 : _GEN_13037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13039 = 7'h45 == _myNewVec_27_T_3[6:0] ? myVec_69 : _GEN_13038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13040 = 7'h46 == _myNewVec_27_T_3[6:0] ? myVec_70 : _GEN_13039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13041 = 7'h47 == _myNewVec_27_T_3[6:0] ? myVec_71 : _GEN_13040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13042 = 7'h48 == _myNewVec_27_T_3[6:0] ? myVec_72 : _GEN_13041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13043 = 7'h49 == _myNewVec_27_T_3[6:0] ? myVec_73 : _GEN_13042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13044 = 7'h4a == _myNewVec_27_T_3[6:0] ? myVec_74 : _GEN_13043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13045 = 7'h4b == _myNewVec_27_T_3[6:0] ? myVec_75 : _GEN_13044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13046 = 7'h4c == _myNewVec_27_T_3[6:0] ? myVec_76 : _GEN_13045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13047 = 7'h4d == _myNewVec_27_T_3[6:0] ? myVec_77 : _GEN_13046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13048 = 7'h4e == _myNewVec_27_T_3[6:0] ? myVec_78 : _GEN_13047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13049 = 7'h4f == _myNewVec_27_T_3[6:0] ? myVec_79 : _GEN_13048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13050 = 7'h50 == _myNewVec_27_T_3[6:0] ? myVec_80 : _GEN_13049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13051 = 7'h51 == _myNewVec_27_T_3[6:0] ? myVec_81 : _GEN_13050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13052 = 7'h52 == _myNewVec_27_T_3[6:0] ? myVec_82 : _GEN_13051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13053 = 7'h53 == _myNewVec_27_T_3[6:0] ? myVec_83 : _GEN_13052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13054 = 7'h54 == _myNewVec_27_T_3[6:0] ? myVec_84 : _GEN_13053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13055 = 7'h55 == _myNewVec_27_T_3[6:0] ? myVec_85 : _GEN_13054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13056 = 7'h56 == _myNewVec_27_T_3[6:0] ? myVec_86 : _GEN_13055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13057 = 7'h57 == _myNewVec_27_T_3[6:0] ? myVec_87 : _GEN_13056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13058 = 7'h58 == _myNewVec_27_T_3[6:0] ? myVec_88 : _GEN_13057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13059 = 7'h59 == _myNewVec_27_T_3[6:0] ? myVec_89 : _GEN_13058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13060 = 7'h5a == _myNewVec_27_T_3[6:0] ? myVec_90 : _GEN_13059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13061 = 7'h5b == _myNewVec_27_T_3[6:0] ? myVec_91 : _GEN_13060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13062 = 7'h5c == _myNewVec_27_T_3[6:0] ? myVec_92 : _GEN_13061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13063 = 7'h5d == _myNewVec_27_T_3[6:0] ? myVec_93 : _GEN_13062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13064 = 7'h5e == _myNewVec_27_T_3[6:0] ? myVec_94 : _GEN_13063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13065 = 7'h5f == _myNewVec_27_T_3[6:0] ? myVec_95 : _GEN_13064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13066 = 7'h60 == _myNewVec_27_T_3[6:0] ? myVec_96 : _GEN_13065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13067 = 7'h61 == _myNewVec_27_T_3[6:0] ? myVec_97 : _GEN_13066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13068 = 7'h62 == _myNewVec_27_T_3[6:0] ? myVec_98 : _GEN_13067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13069 = 7'h63 == _myNewVec_27_T_3[6:0] ? myVec_99 : _GEN_13068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13070 = 7'h64 == _myNewVec_27_T_3[6:0] ? myVec_100 : _GEN_13069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13071 = 7'h65 == _myNewVec_27_T_3[6:0] ? myVec_101 : _GEN_13070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13072 = 7'h66 == _myNewVec_27_T_3[6:0] ? myVec_102 : _GEN_13071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13073 = 7'h67 == _myNewVec_27_T_3[6:0] ? myVec_103 : _GEN_13072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13074 = 7'h68 == _myNewVec_27_T_3[6:0] ? myVec_104 : _GEN_13073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13075 = 7'h69 == _myNewVec_27_T_3[6:0] ? myVec_105 : _GEN_13074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13076 = 7'h6a == _myNewVec_27_T_3[6:0] ? myVec_106 : _GEN_13075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13077 = 7'h6b == _myNewVec_27_T_3[6:0] ? myVec_107 : _GEN_13076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13078 = 7'h6c == _myNewVec_27_T_3[6:0] ? myVec_108 : _GEN_13077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13079 = 7'h6d == _myNewVec_27_T_3[6:0] ? myVec_109 : _GEN_13078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13080 = 7'h6e == _myNewVec_27_T_3[6:0] ? myVec_110 : _GEN_13079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13081 = 7'h6f == _myNewVec_27_T_3[6:0] ? myVec_111 : _GEN_13080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13082 = 7'h70 == _myNewVec_27_T_3[6:0] ? myVec_112 : _GEN_13081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13083 = 7'h71 == _myNewVec_27_T_3[6:0] ? myVec_113 : _GEN_13082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13084 = 7'h72 == _myNewVec_27_T_3[6:0] ? myVec_114 : _GEN_13083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13085 = 7'h73 == _myNewVec_27_T_3[6:0] ? myVec_115 : _GEN_13084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13086 = 7'h74 == _myNewVec_27_T_3[6:0] ? myVec_116 : _GEN_13085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13087 = 7'h75 == _myNewVec_27_T_3[6:0] ? myVec_117 : _GEN_13086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13088 = 7'h76 == _myNewVec_27_T_3[6:0] ? myVec_118 : _GEN_13087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13089 = 7'h77 == _myNewVec_27_T_3[6:0] ? myVec_119 : _GEN_13088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13090 = 7'h78 == _myNewVec_27_T_3[6:0] ? myVec_120 : _GEN_13089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13091 = 7'h79 == _myNewVec_27_T_3[6:0] ? myVec_121 : _GEN_13090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13092 = 7'h7a == _myNewVec_27_T_3[6:0] ? myVec_122 : _GEN_13091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13093 = 7'h7b == _myNewVec_27_T_3[6:0] ? myVec_123 : _GEN_13092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13094 = 7'h7c == _myNewVec_27_T_3[6:0] ? myVec_124 : _GEN_13093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13095 = 7'h7d == _myNewVec_27_T_3[6:0] ? myVec_125 : _GEN_13094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13096 = 7'h7e == _myNewVec_27_T_3[6:0] ? myVec_126 : _GEN_13095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_27 = 7'h7f == _myNewVec_27_T_3[6:0] ? myVec_127 : _GEN_13096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_26_T_3 = _myNewVec_127_T_1 + 16'h65; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_13099 = 7'h1 == _myNewVec_26_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13100 = 7'h2 == _myNewVec_26_T_3[6:0] ? myVec_2 : _GEN_13099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13101 = 7'h3 == _myNewVec_26_T_3[6:0] ? myVec_3 : _GEN_13100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13102 = 7'h4 == _myNewVec_26_T_3[6:0] ? myVec_4 : _GEN_13101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13103 = 7'h5 == _myNewVec_26_T_3[6:0] ? myVec_5 : _GEN_13102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13104 = 7'h6 == _myNewVec_26_T_3[6:0] ? myVec_6 : _GEN_13103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13105 = 7'h7 == _myNewVec_26_T_3[6:0] ? myVec_7 : _GEN_13104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13106 = 7'h8 == _myNewVec_26_T_3[6:0] ? myVec_8 : _GEN_13105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13107 = 7'h9 == _myNewVec_26_T_3[6:0] ? myVec_9 : _GEN_13106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13108 = 7'ha == _myNewVec_26_T_3[6:0] ? myVec_10 : _GEN_13107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13109 = 7'hb == _myNewVec_26_T_3[6:0] ? myVec_11 : _GEN_13108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13110 = 7'hc == _myNewVec_26_T_3[6:0] ? myVec_12 : _GEN_13109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13111 = 7'hd == _myNewVec_26_T_3[6:0] ? myVec_13 : _GEN_13110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13112 = 7'he == _myNewVec_26_T_3[6:0] ? myVec_14 : _GEN_13111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13113 = 7'hf == _myNewVec_26_T_3[6:0] ? myVec_15 : _GEN_13112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13114 = 7'h10 == _myNewVec_26_T_3[6:0] ? myVec_16 : _GEN_13113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13115 = 7'h11 == _myNewVec_26_T_3[6:0] ? myVec_17 : _GEN_13114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13116 = 7'h12 == _myNewVec_26_T_3[6:0] ? myVec_18 : _GEN_13115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13117 = 7'h13 == _myNewVec_26_T_3[6:0] ? myVec_19 : _GEN_13116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13118 = 7'h14 == _myNewVec_26_T_3[6:0] ? myVec_20 : _GEN_13117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13119 = 7'h15 == _myNewVec_26_T_3[6:0] ? myVec_21 : _GEN_13118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13120 = 7'h16 == _myNewVec_26_T_3[6:0] ? myVec_22 : _GEN_13119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13121 = 7'h17 == _myNewVec_26_T_3[6:0] ? myVec_23 : _GEN_13120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13122 = 7'h18 == _myNewVec_26_T_3[6:0] ? myVec_24 : _GEN_13121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13123 = 7'h19 == _myNewVec_26_T_3[6:0] ? myVec_25 : _GEN_13122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13124 = 7'h1a == _myNewVec_26_T_3[6:0] ? myVec_26 : _GEN_13123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13125 = 7'h1b == _myNewVec_26_T_3[6:0] ? myVec_27 : _GEN_13124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13126 = 7'h1c == _myNewVec_26_T_3[6:0] ? myVec_28 : _GEN_13125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13127 = 7'h1d == _myNewVec_26_T_3[6:0] ? myVec_29 : _GEN_13126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13128 = 7'h1e == _myNewVec_26_T_3[6:0] ? myVec_30 : _GEN_13127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13129 = 7'h1f == _myNewVec_26_T_3[6:0] ? myVec_31 : _GEN_13128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13130 = 7'h20 == _myNewVec_26_T_3[6:0] ? myVec_32 : _GEN_13129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13131 = 7'h21 == _myNewVec_26_T_3[6:0] ? myVec_33 : _GEN_13130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13132 = 7'h22 == _myNewVec_26_T_3[6:0] ? myVec_34 : _GEN_13131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13133 = 7'h23 == _myNewVec_26_T_3[6:0] ? myVec_35 : _GEN_13132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13134 = 7'h24 == _myNewVec_26_T_3[6:0] ? myVec_36 : _GEN_13133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13135 = 7'h25 == _myNewVec_26_T_3[6:0] ? myVec_37 : _GEN_13134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13136 = 7'h26 == _myNewVec_26_T_3[6:0] ? myVec_38 : _GEN_13135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13137 = 7'h27 == _myNewVec_26_T_3[6:0] ? myVec_39 : _GEN_13136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13138 = 7'h28 == _myNewVec_26_T_3[6:0] ? myVec_40 : _GEN_13137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13139 = 7'h29 == _myNewVec_26_T_3[6:0] ? myVec_41 : _GEN_13138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13140 = 7'h2a == _myNewVec_26_T_3[6:0] ? myVec_42 : _GEN_13139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13141 = 7'h2b == _myNewVec_26_T_3[6:0] ? myVec_43 : _GEN_13140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13142 = 7'h2c == _myNewVec_26_T_3[6:0] ? myVec_44 : _GEN_13141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13143 = 7'h2d == _myNewVec_26_T_3[6:0] ? myVec_45 : _GEN_13142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13144 = 7'h2e == _myNewVec_26_T_3[6:0] ? myVec_46 : _GEN_13143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13145 = 7'h2f == _myNewVec_26_T_3[6:0] ? myVec_47 : _GEN_13144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13146 = 7'h30 == _myNewVec_26_T_3[6:0] ? myVec_48 : _GEN_13145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13147 = 7'h31 == _myNewVec_26_T_3[6:0] ? myVec_49 : _GEN_13146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13148 = 7'h32 == _myNewVec_26_T_3[6:0] ? myVec_50 : _GEN_13147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13149 = 7'h33 == _myNewVec_26_T_3[6:0] ? myVec_51 : _GEN_13148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13150 = 7'h34 == _myNewVec_26_T_3[6:0] ? myVec_52 : _GEN_13149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13151 = 7'h35 == _myNewVec_26_T_3[6:0] ? myVec_53 : _GEN_13150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13152 = 7'h36 == _myNewVec_26_T_3[6:0] ? myVec_54 : _GEN_13151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13153 = 7'h37 == _myNewVec_26_T_3[6:0] ? myVec_55 : _GEN_13152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13154 = 7'h38 == _myNewVec_26_T_3[6:0] ? myVec_56 : _GEN_13153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13155 = 7'h39 == _myNewVec_26_T_3[6:0] ? myVec_57 : _GEN_13154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13156 = 7'h3a == _myNewVec_26_T_3[6:0] ? myVec_58 : _GEN_13155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13157 = 7'h3b == _myNewVec_26_T_3[6:0] ? myVec_59 : _GEN_13156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13158 = 7'h3c == _myNewVec_26_T_3[6:0] ? myVec_60 : _GEN_13157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13159 = 7'h3d == _myNewVec_26_T_3[6:0] ? myVec_61 : _GEN_13158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13160 = 7'h3e == _myNewVec_26_T_3[6:0] ? myVec_62 : _GEN_13159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13161 = 7'h3f == _myNewVec_26_T_3[6:0] ? myVec_63 : _GEN_13160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13162 = 7'h40 == _myNewVec_26_T_3[6:0] ? myVec_64 : _GEN_13161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13163 = 7'h41 == _myNewVec_26_T_3[6:0] ? myVec_65 : _GEN_13162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13164 = 7'h42 == _myNewVec_26_T_3[6:0] ? myVec_66 : _GEN_13163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13165 = 7'h43 == _myNewVec_26_T_3[6:0] ? myVec_67 : _GEN_13164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13166 = 7'h44 == _myNewVec_26_T_3[6:0] ? myVec_68 : _GEN_13165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13167 = 7'h45 == _myNewVec_26_T_3[6:0] ? myVec_69 : _GEN_13166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13168 = 7'h46 == _myNewVec_26_T_3[6:0] ? myVec_70 : _GEN_13167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13169 = 7'h47 == _myNewVec_26_T_3[6:0] ? myVec_71 : _GEN_13168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13170 = 7'h48 == _myNewVec_26_T_3[6:0] ? myVec_72 : _GEN_13169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13171 = 7'h49 == _myNewVec_26_T_3[6:0] ? myVec_73 : _GEN_13170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13172 = 7'h4a == _myNewVec_26_T_3[6:0] ? myVec_74 : _GEN_13171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13173 = 7'h4b == _myNewVec_26_T_3[6:0] ? myVec_75 : _GEN_13172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13174 = 7'h4c == _myNewVec_26_T_3[6:0] ? myVec_76 : _GEN_13173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13175 = 7'h4d == _myNewVec_26_T_3[6:0] ? myVec_77 : _GEN_13174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13176 = 7'h4e == _myNewVec_26_T_3[6:0] ? myVec_78 : _GEN_13175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13177 = 7'h4f == _myNewVec_26_T_3[6:0] ? myVec_79 : _GEN_13176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13178 = 7'h50 == _myNewVec_26_T_3[6:0] ? myVec_80 : _GEN_13177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13179 = 7'h51 == _myNewVec_26_T_3[6:0] ? myVec_81 : _GEN_13178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13180 = 7'h52 == _myNewVec_26_T_3[6:0] ? myVec_82 : _GEN_13179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13181 = 7'h53 == _myNewVec_26_T_3[6:0] ? myVec_83 : _GEN_13180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13182 = 7'h54 == _myNewVec_26_T_3[6:0] ? myVec_84 : _GEN_13181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13183 = 7'h55 == _myNewVec_26_T_3[6:0] ? myVec_85 : _GEN_13182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13184 = 7'h56 == _myNewVec_26_T_3[6:0] ? myVec_86 : _GEN_13183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13185 = 7'h57 == _myNewVec_26_T_3[6:0] ? myVec_87 : _GEN_13184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13186 = 7'h58 == _myNewVec_26_T_3[6:0] ? myVec_88 : _GEN_13185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13187 = 7'h59 == _myNewVec_26_T_3[6:0] ? myVec_89 : _GEN_13186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13188 = 7'h5a == _myNewVec_26_T_3[6:0] ? myVec_90 : _GEN_13187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13189 = 7'h5b == _myNewVec_26_T_3[6:0] ? myVec_91 : _GEN_13188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13190 = 7'h5c == _myNewVec_26_T_3[6:0] ? myVec_92 : _GEN_13189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13191 = 7'h5d == _myNewVec_26_T_3[6:0] ? myVec_93 : _GEN_13190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13192 = 7'h5e == _myNewVec_26_T_3[6:0] ? myVec_94 : _GEN_13191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13193 = 7'h5f == _myNewVec_26_T_3[6:0] ? myVec_95 : _GEN_13192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13194 = 7'h60 == _myNewVec_26_T_3[6:0] ? myVec_96 : _GEN_13193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13195 = 7'h61 == _myNewVec_26_T_3[6:0] ? myVec_97 : _GEN_13194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13196 = 7'h62 == _myNewVec_26_T_3[6:0] ? myVec_98 : _GEN_13195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13197 = 7'h63 == _myNewVec_26_T_3[6:0] ? myVec_99 : _GEN_13196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13198 = 7'h64 == _myNewVec_26_T_3[6:0] ? myVec_100 : _GEN_13197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13199 = 7'h65 == _myNewVec_26_T_3[6:0] ? myVec_101 : _GEN_13198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13200 = 7'h66 == _myNewVec_26_T_3[6:0] ? myVec_102 : _GEN_13199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13201 = 7'h67 == _myNewVec_26_T_3[6:0] ? myVec_103 : _GEN_13200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13202 = 7'h68 == _myNewVec_26_T_3[6:0] ? myVec_104 : _GEN_13201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13203 = 7'h69 == _myNewVec_26_T_3[6:0] ? myVec_105 : _GEN_13202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13204 = 7'h6a == _myNewVec_26_T_3[6:0] ? myVec_106 : _GEN_13203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13205 = 7'h6b == _myNewVec_26_T_3[6:0] ? myVec_107 : _GEN_13204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13206 = 7'h6c == _myNewVec_26_T_3[6:0] ? myVec_108 : _GEN_13205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13207 = 7'h6d == _myNewVec_26_T_3[6:0] ? myVec_109 : _GEN_13206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13208 = 7'h6e == _myNewVec_26_T_3[6:0] ? myVec_110 : _GEN_13207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13209 = 7'h6f == _myNewVec_26_T_3[6:0] ? myVec_111 : _GEN_13208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13210 = 7'h70 == _myNewVec_26_T_3[6:0] ? myVec_112 : _GEN_13209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13211 = 7'h71 == _myNewVec_26_T_3[6:0] ? myVec_113 : _GEN_13210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13212 = 7'h72 == _myNewVec_26_T_3[6:0] ? myVec_114 : _GEN_13211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13213 = 7'h73 == _myNewVec_26_T_3[6:0] ? myVec_115 : _GEN_13212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13214 = 7'h74 == _myNewVec_26_T_3[6:0] ? myVec_116 : _GEN_13213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13215 = 7'h75 == _myNewVec_26_T_3[6:0] ? myVec_117 : _GEN_13214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13216 = 7'h76 == _myNewVec_26_T_3[6:0] ? myVec_118 : _GEN_13215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13217 = 7'h77 == _myNewVec_26_T_3[6:0] ? myVec_119 : _GEN_13216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13218 = 7'h78 == _myNewVec_26_T_3[6:0] ? myVec_120 : _GEN_13217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13219 = 7'h79 == _myNewVec_26_T_3[6:0] ? myVec_121 : _GEN_13218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13220 = 7'h7a == _myNewVec_26_T_3[6:0] ? myVec_122 : _GEN_13219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13221 = 7'h7b == _myNewVec_26_T_3[6:0] ? myVec_123 : _GEN_13220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13222 = 7'h7c == _myNewVec_26_T_3[6:0] ? myVec_124 : _GEN_13221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13223 = 7'h7d == _myNewVec_26_T_3[6:0] ? myVec_125 : _GEN_13222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13224 = 7'h7e == _myNewVec_26_T_3[6:0] ? myVec_126 : _GEN_13223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_26 = 7'h7f == _myNewVec_26_T_3[6:0] ? myVec_127 : _GEN_13224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_25_T_3 = _myNewVec_127_T_1 + 16'h66; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_13227 = 7'h1 == _myNewVec_25_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13228 = 7'h2 == _myNewVec_25_T_3[6:0] ? myVec_2 : _GEN_13227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13229 = 7'h3 == _myNewVec_25_T_3[6:0] ? myVec_3 : _GEN_13228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13230 = 7'h4 == _myNewVec_25_T_3[6:0] ? myVec_4 : _GEN_13229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13231 = 7'h5 == _myNewVec_25_T_3[6:0] ? myVec_5 : _GEN_13230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13232 = 7'h6 == _myNewVec_25_T_3[6:0] ? myVec_6 : _GEN_13231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13233 = 7'h7 == _myNewVec_25_T_3[6:0] ? myVec_7 : _GEN_13232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13234 = 7'h8 == _myNewVec_25_T_3[6:0] ? myVec_8 : _GEN_13233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13235 = 7'h9 == _myNewVec_25_T_3[6:0] ? myVec_9 : _GEN_13234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13236 = 7'ha == _myNewVec_25_T_3[6:0] ? myVec_10 : _GEN_13235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13237 = 7'hb == _myNewVec_25_T_3[6:0] ? myVec_11 : _GEN_13236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13238 = 7'hc == _myNewVec_25_T_3[6:0] ? myVec_12 : _GEN_13237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13239 = 7'hd == _myNewVec_25_T_3[6:0] ? myVec_13 : _GEN_13238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13240 = 7'he == _myNewVec_25_T_3[6:0] ? myVec_14 : _GEN_13239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13241 = 7'hf == _myNewVec_25_T_3[6:0] ? myVec_15 : _GEN_13240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13242 = 7'h10 == _myNewVec_25_T_3[6:0] ? myVec_16 : _GEN_13241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13243 = 7'h11 == _myNewVec_25_T_3[6:0] ? myVec_17 : _GEN_13242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13244 = 7'h12 == _myNewVec_25_T_3[6:0] ? myVec_18 : _GEN_13243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13245 = 7'h13 == _myNewVec_25_T_3[6:0] ? myVec_19 : _GEN_13244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13246 = 7'h14 == _myNewVec_25_T_3[6:0] ? myVec_20 : _GEN_13245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13247 = 7'h15 == _myNewVec_25_T_3[6:0] ? myVec_21 : _GEN_13246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13248 = 7'h16 == _myNewVec_25_T_3[6:0] ? myVec_22 : _GEN_13247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13249 = 7'h17 == _myNewVec_25_T_3[6:0] ? myVec_23 : _GEN_13248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13250 = 7'h18 == _myNewVec_25_T_3[6:0] ? myVec_24 : _GEN_13249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13251 = 7'h19 == _myNewVec_25_T_3[6:0] ? myVec_25 : _GEN_13250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13252 = 7'h1a == _myNewVec_25_T_3[6:0] ? myVec_26 : _GEN_13251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13253 = 7'h1b == _myNewVec_25_T_3[6:0] ? myVec_27 : _GEN_13252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13254 = 7'h1c == _myNewVec_25_T_3[6:0] ? myVec_28 : _GEN_13253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13255 = 7'h1d == _myNewVec_25_T_3[6:0] ? myVec_29 : _GEN_13254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13256 = 7'h1e == _myNewVec_25_T_3[6:0] ? myVec_30 : _GEN_13255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13257 = 7'h1f == _myNewVec_25_T_3[6:0] ? myVec_31 : _GEN_13256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13258 = 7'h20 == _myNewVec_25_T_3[6:0] ? myVec_32 : _GEN_13257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13259 = 7'h21 == _myNewVec_25_T_3[6:0] ? myVec_33 : _GEN_13258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13260 = 7'h22 == _myNewVec_25_T_3[6:0] ? myVec_34 : _GEN_13259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13261 = 7'h23 == _myNewVec_25_T_3[6:0] ? myVec_35 : _GEN_13260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13262 = 7'h24 == _myNewVec_25_T_3[6:0] ? myVec_36 : _GEN_13261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13263 = 7'h25 == _myNewVec_25_T_3[6:0] ? myVec_37 : _GEN_13262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13264 = 7'h26 == _myNewVec_25_T_3[6:0] ? myVec_38 : _GEN_13263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13265 = 7'h27 == _myNewVec_25_T_3[6:0] ? myVec_39 : _GEN_13264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13266 = 7'h28 == _myNewVec_25_T_3[6:0] ? myVec_40 : _GEN_13265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13267 = 7'h29 == _myNewVec_25_T_3[6:0] ? myVec_41 : _GEN_13266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13268 = 7'h2a == _myNewVec_25_T_3[6:0] ? myVec_42 : _GEN_13267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13269 = 7'h2b == _myNewVec_25_T_3[6:0] ? myVec_43 : _GEN_13268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13270 = 7'h2c == _myNewVec_25_T_3[6:0] ? myVec_44 : _GEN_13269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13271 = 7'h2d == _myNewVec_25_T_3[6:0] ? myVec_45 : _GEN_13270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13272 = 7'h2e == _myNewVec_25_T_3[6:0] ? myVec_46 : _GEN_13271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13273 = 7'h2f == _myNewVec_25_T_3[6:0] ? myVec_47 : _GEN_13272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13274 = 7'h30 == _myNewVec_25_T_3[6:0] ? myVec_48 : _GEN_13273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13275 = 7'h31 == _myNewVec_25_T_3[6:0] ? myVec_49 : _GEN_13274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13276 = 7'h32 == _myNewVec_25_T_3[6:0] ? myVec_50 : _GEN_13275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13277 = 7'h33 == _myNewVec_25_T_3[6:0] ? myVec_51 : _GEN_13276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13278 = 7'h34 == _myNewVec_25_T_3[6:0] ? myVec_52 : _GEN_13277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13279 = 7'h35 == _myNewVec_25_T_3[6:0] ? myVec_53 : _GEN_13278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13280 = 7'h36 == _myNewVec_25_T_3[6:0] ? myVec_54 : _GEN_13279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13281 = 7'h37 == _myNewVec_25_T_3[6:0] ? myVec_55 : _GEN_13280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13282 = 7'h38 == _myNewVec_25_T_3[6:0] ? myVec_56 : _GEN_13281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13283 = 7'h39 == _myNewVec_25_T_3[6:0] ? myVec_57 : _GEN_13282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13284 = 7'h3a == _myNewVec_25_T_3[6:0] ? myVec_58 : _GEN_13283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13285 = 7'h3b == _myNewVec_25_T_3[6:0] ? myVec_59 : _GEN_13284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13286 = 7'h3c == _myNewVec_25_T_3[6:0] ? myVec_60 : _GEN_13285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13287 = 7'h3d == _myNewVec_25_T_3[6:0] ? myVec_61 : _GEN_13286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13288 = 7'h3e == _myNewVec_25_T_3[6:0] ? myVec_62 : _GEN_13287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13289 = 7'h3f == _myNewVec_25_T_3[6:0] ? myVec_63 : _GEN_13288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13290 = 7'h40 == _myNewVec_25_T_3[6:0] ? myVec_64 : _GEN_13289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13291 = 7'h41 == _myNewVec_25_T_3[6:0] ? myVec_65 : _GEN_13290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13292 = 7'h42 == _myNewVec_25_T_3[6:0] ? myVec_66 : _GEN_13291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13293 = 7'h43 == _myNewVec_25_T_3[6:0] ? myVec_67 : _GEN_13292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13294 = 7'h44 == _myNewVec_25_T_3[6:0] ? myVec_68 : _GEN_13293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13295 = 7'h45 == _myNewVec_25_T_3[6:0] ? myVec_69 : _GEN_13294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13296 = 7'h46 == _myNewVec_25_T_3[6:0] ? myVec_70 : _GEN_13295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13297 = 7'h47 == _myNewVec_25_T_3[6:0] ? myVec_71 : _GEN_13296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13298 = 7'h48 == _myNewVec_25_T_3[6:0] ? myVec_72 : _GEN_13297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13299 = 7'h49 == _myNewVec_25_T_3[6:0] ? myVec_73 : _GEN_13298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13300 = 7'h4a == _myNewVec_25_T_3[6:0] ? myVec_74 : _GEN_13299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13301 = 7'h4b == _myNewVec_25_T_3[6:0] ? myVec_75 : _GEN_13300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13302 = 7'h4c == _myNewVec_25_T_3[6:0] ? myVec_76 : _GEN_13301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13303 = 7'h4d == _myNewVec_25_T_3[6:0] ? myVec_77 : _GEN_13302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13304 = 7'h4e == _myNewVec_25_T_3[6:0] ? myVec_78 : _GEN_13303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13305 = 7'h4f == _myNewVec_25_T_3[6:0] ? myVec_79 : _GEN_13304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13306 = 7'h50 == _myNewVec_25_T_3[6:0] ? myVec_80 : _GEN_13305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13307 = 7'h51 == _myNewVec_25_T_3[6:0] ? myVec_81 : _GEN_13306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13308 = 7'h52 == _myNewVec_25_T_3[6:0] ? myVec_82 : _GEN_13307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13309 = 7'h53 == _myNewVec_25_T_3[6:0] ? myVec_83 : _GEN_13308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13310 = 7'h54 == _myNewVec_25_T_3[6:0] ? myVec_84 : _GEN_13309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13311 = 7'h55 == _myNewVec_25_T_3[6:0] ? myVec_85 : _GEN_13310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13312 = 7'h56 == _myNewVec_25_T_3[6:0] ? myVec_86 : _GEN_13311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13313 = 7'h57 == _myNewVec_25_T_3[6:0] ? myVec_87 : _GEN_13312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13314 = 7'h58 == _myNewVec_25_T_3[6:0] ? myVec_88 : _GEN_13313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13315 = 7'h59 == _myNewVec_25_T_3[6:0] ? myVec_89 : _GEN_13314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13316 = 7'h5a == _myNewVec_25_T_3[6:0] ? myVec_90 : _GEN_13315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13317 = 7'h5b == _myNewVec_25_T_3[6:0] ? myVec_91 : _GEN_13316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13318 = 7'h5c == _myNewVec_25_T_3[6:0] ? myVec_92 : _GEN_13317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13319 = 7'h5d == _myNewVec_25_T_3[6:0] ? myVec_93 : _GEN_13318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13320 = 7'h5e == _myNewVec_25_T_3[6:0] ? myVec_94 : _GEN_13319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13321 = 7'h5f == _myNewVec_25_T_3[6:0] ? myVec_95 : _GEN_13320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13322 = 7'h60 == _myNewVec_25_T_3[6:0] ? myVec_96 : _GEN_13321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13323 = 7'h61 == _myNewVec_25_T_3[6:0] ? myVec_97 : _GEN_13322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13324 = 7'h62 == _myNewVec_25_T_3[6:0] ? myVec_98 : _GEN_13323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13325 = 7'h63 == _myNewVec_25_T_3[6:0] ? myVec_99 : _GEN_13324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13326 = 7'h64 == _myNewVec_25_T_3[6:0] ? myVec_100 : _GEN_13325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13327 = 7'h65 == _myNewVec_25_T_3[6:0] ? myVec_101 : _GEN_13326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13328 = 7'h66 == _myNewVec_25_T_3[6:0] ? myVec_102 : _GEN_13327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13329 = 7'h67 == _myNewVec_25_T_3[6:0] ? myVec_103 : _GEN_13328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13330 = 7'h68 == _myNewVec_25_T_3[6:0] ? myVec_104 : _GEN_13329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13331 = 7'h69 == _myNewVec_25_T_3[6:0] ? myVec_105 : _GEN_13330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13332 = 7'h6a == _myNewVec_25_T_3[6:0] ? myVec_106 : _GEN_13331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13333 = 7'h6b == _myNewVec_25_T_3[6:0] ? myVec_107 : _GEN_13332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13334 = 7'h6c == _myNewVec_25_T_3[6:0] ? myVec_108 : _GEN_13333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13335 = 7'h6d == _myNewVec_25_T_3[6:0] ? myVec_109 : _GEN_13334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13336 = 7'h6e == _myNewVec_25_T_3[6:0] ? myVec_110 : _GEN_13335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13337 = 7'h6f == _myNewVec_25_T_3[6:0] ? myVec_111 : _GEN_13336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13338 = 7'h70 == _myNewVec_25_T_3[6:0] ? myVec_112 : _GEN_13337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13339 = 7'h71 == _myNewVec_25_T_3[6:0] ? myVec_113 : _GEN_13338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13340 = 7'h72 == _myNewVec_25_T_3[6:0] ? myVec_114 : _GEN_13339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13341 = 7'h73 == _myNewVec_25_T_3[6:0] ? myVec_115 : _GEN_13340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13342 = 7'h74 == _myNewVec_25_T_3[6:0] ? myVec_116 : _GEN_13341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13343 = 7'h75 == _myNewVec_25_T_3[6:0] ? myVec_117 : _GEN_13342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13344 = 7'h76 == _myNewVec_25_T_3[6:0] ? myVec_118 : _GEN_13343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13345 = 7'h77 == _myNewVec_25_T_3[6:0] ? myVec_119 : _GEN_13344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13346 = 7'h78 == _myNewVec_25_T_3[6:0] ? myVec_120 : _GEN_13345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13347 = 7'h79 == _myNewVec_25_T_3[6:0] ? myVec_121 : _GEN_13346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13348 = 7'h7a == _myNewVec_25_T_3[6:0] ? myVec_122 : _GEN_13347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13349 = 7'h7b == _myNewVec_25_T_3[6:0] ? myVec_123 : _GEN_13348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13350 = 7'h7c == _myNewVec_25_T_3[6:0] ? myVec_124 : _GEN_13349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13351 = 7'h7d == _myNewVec_25_T_3[6:0] ? myVec_125 : _GEN_13350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13352 = 7'h7e == _myNewVec_25_T_3[6:0] ? myVec_126 : _GEN_13351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_25 = 7'h7f == _myNewVec_25_T_3[6:0] ? myVec_127 : _GEN_13352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_24_T_3 = _myNewVec_127_T_1 + 16'h67; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_13355 = 7'h1 == _myNewVec_24_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13356 = 7'h2 == _myNewVec_24_T_3[6:0] ? myVec_2 : _GEN_13355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13357 = 7'h3 == _myNewVec_24_T_3[6:0] ? myVec_3 : _GEN_13356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13358 = 7'h4 == _myNewVec_24_T_3[6:0] ? myVec_4 : _GEN_13357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13359 = 7'h5 == _myNewVec_24_T_3[6:0] ? myVec_5 : _GEN_13358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13360 = 7'h6 == _myNewVec_24_T_3[6:0] ? myVec_6 : _GEN_13359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13361 = 7'h7 == _myNewVec_24_T_3[6:0] ? myVec_7 : _GEN_13360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13362 = 7'h8 == _myNewVec_24_T_3[6:0] ? myVec_8 : _GEN_13361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13363 = 7'h9 == _myNewVec_24_T_3[6:0] ? myVec_9 : _GEN_13362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13364 = 7'ha == _myNewVec_24_T_3[6:0] ? myVec_10 : _GEN_13363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13365 = 7'hb == _myNewVec_24_T_3[6:0] ? myVec_11 : _GEN_13364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13366 = 7'hc == _myNewVec_24_T_3[6:0] ? myVec_12 : _GEN_13365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13367 = 7'hd == _myNewVec_24_T_3[6:0] ? myVec_13 : _GEN_13366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13368 = 7'he == _myNewVec_24_T_3[6:0] ? myVec_14 : _GEN_13367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13369 = 7'hf == _myNewVec_24_T_3[6:0] ? myVec_15 : _GEN_13368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13370 = 7'h10 == _myNewVec_24_T_3[6:0] ? myVec_16 : _GEN_13369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13371 = 7'h11 == _myNewVec_24_T_3[6:0] ? myVec_17 : _GEN_13370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13372 = 7'h12 == _myNewVec_24_T_3[6:0] ? myVec_18 : _GEN_13371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13373 = 7'h13 == _myNewVec_24_T_3[6:0] ? myVec_19 : _GEN_13372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13374 = 7'h14 == _myNewVec_24_T_3[6:0] ? myVec_20 : _GEN_13373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13375 = 7'h15 == _myNewVec_24_T_3[6:0] ? myVec_21 : _GEN_13374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13376 = 7'h16 == _myNewVec_24_T_3[6:0] ? myVec_22 : _GEN_13375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13377 = 7'h17 == _myNewVec_24_T_3[6:0] ? myVec_23 : _GEN_13376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13378 = 7'h18 == _myNewVec_24_T_3[6:0] ? myVec_24 : _GEN_13377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13379 = 7'h19 == _myNewVec_24_T_3[6:0] ? myVec_25 : _GEN_13378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13380 = 7'h1a == _myNewVec_24_T_3[6:0] ? myVec_26 : _GEN_13379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13381 = 7'h1b == _myNewVec_24_T_3[6:0] ? myVec_27 : _GEN_13380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13382 = 7'h1c == _myNewVec_24_T_3[6:0] ? myVec_28 : _GEN_13381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13383 = 7'h1d == _myNewVec_24_T_3[6:0] ? myVec_29 : _GEN_13382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13384 = 7'h1e == _myNewVec_24_T_3[6:0] ? myVec_30 : _GEN_13383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13385 = 7'h1f == _myNewVec_24_T_3[6:0] ? myVec_31 : _GEN_13384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13386 = 7'h20 == _myNewVec_24_T_3[6:0] ? myVec_32 : _GEN_13385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13387 = 7'h21 == _myNewVec_24_T_3[6:0] ? myVec_33 : _GEN_13386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13388 = 7'h22 == _myNewVec_24_T_3[6:0] ? myVec_34 : _GEN_13387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13389 = 7'h23 == _myNewVec_24_T_3[6:0] ? myVec_35 : _GEN_13388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13390 = 7'h24 == _myNewVec_24_T_3[6:0] ? myVec_36 : _GEN_13389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13391 = 7'h25 == _myNewVec_24_T_3[6:0] ? myVec_37 : _GEN_13390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13392 = 7'h26 == _myNewVec_24_T_3[6:0] ? myVec_38 : _GEN_13391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13393 = 7'h27 == _myNewVec_24_T_3[6:0] ? myVec_39 : _GEN_13392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13394 = 7'h28 == _myNewVec_24_T_3[6:0] ? myVec_40 : _GEN_13393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13395 = 7'h29 == _myNewVec_24_T_3[6:0] ? myVec_41 : _GEN_13394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13396 = 7'h2a == _myNewVec_24_T_3[6:0] ? myVec_42 : _GEN_13395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13397 = 7'h2b == _myNewVec_24_T_3[6:0] ? myVec_43 : _GEN_13396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13398 = 7'h2c == _myNewVec_24_T_3[6:0] ? myVec_44 : _GEN_13397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13399 = 7'h2d == _myNewVec_24_T_3[6:0] ? myVec_45 : _GEN_13398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13400 = 7'h2e == _myNewVec_24_T_3[6:0] ? myVec_46 : _GEN_13399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13401 = 7'h2f == _myNewVec_24_T_3[6:0] ? myVec_47 : _GEN_13400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13402 = 7'h30 == _myNewVec_24_T_3[6:0] ? myVec_48 : _GEN_13401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13403 = 7'h31 == _myNewVec_24_T_3[6:0] ? myVec_49 : _GEN_13402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13404 = 7'h32 == _myNewVec_24_T_3[6:0] ? myVec_50 : _GEN_13403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13405 = 7'h33 == _myNewVec_24_T_3[6:0] ? myVec_51 : _GEN_13404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13406 = 7'h34 == _myNewVec_24_T_3[6:0] ? myVec_52 : _GEN_13405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13407 = 7'h35 == _myNewVec_24_T_3[6:0] ? myVec_53 : _GEN_13406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13408 = 7'h36 == _myNewVec_24_T_3[6:0] ? myVec_54 : _GEN_13407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13409 = 7'h37 == _myNewVec_24_T_3[6:0] ? myVec_55 : _GEN_13408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13410 = 7'h38 == _myNewVec_24_T_3[6:0] ? myVec_56 : _GEN_13409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13411 = 7'h39 == _myNewVec_24_T_3[6:0] ? myVec_57 : _GEN_13410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13412 = 7'h3a == _myNewVec_24_T_3[6:0] ? myVec_58 : _GEN_13411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13413 = 7'h3b == _myNewVec_24_T_3[6:0] ? myVec_59 : _GEN_13412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13414 = 7'h3c == _myNewVec_24_T_3[6:0] ? myVec_60 : _GEN_13413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13415 = 7'h3d == _myNewVec_24_T_3[6:0] ? myVec_61 : _GEN_13414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13416 = 7'h3e == _myNewVec_24_T_3[6:0] ? myVec_62 : _GEN_13415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13417 = 7'h3f == _myNewVec_24_T_3[6:0] ? myVec_63 : _GEN_13416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13418 = 7'h40 == _myNewVec_24_T_3[6:0] ? myVec_64 : _GEN_13417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13419 = 7'h41 == _myNewVec_24_T_3[6:0] ? myVec_65 : _GEN_13418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13420 = 7'h42 == _myNewVec_24_T_3[6:0] ? myVec_66 : _GEN_13419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13421 = 7'h43 == _myNewVec_24_T_3[6:0] ? myVec_67 : _GEN_13420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13422 = 7'h44 == _myNewVec_24_T_3[6:0] ? myVec_68 : _GEN_13421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13423 = 7'h45 == _myNewVec_24_T_3[6:0] ? myVec_69 : _GEN_13422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13424 = 7'h46 == _myNewVec_24_T_3[6:0] ? myVec_70 : _GEN_13423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13425 = 7'h47 == _myNewVec_24_T_3[6:0] ? myVec_71 : _GEN_13424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13426 = 7'h48 == _myNewVec_24_T_3[6:0] ? myVec_72 : _GEN_13425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13427 = 7'h49 == _myNewVec_24_T_3[6:0] ? myVec_73 : _GEN_13426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13428 = 7'h4a == _myNewVec_24_T_3[6:0] ? myVec_74 : _GEN_13427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13429 = 7'h4b == _myNewVec_24_T_3[6:0] ? myVec_75 : _GEN_13428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13430 = 7'h4c == _myNewVec_24_T_3[6:0] ? myVec_76 : _GEN_13429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13431 = 7'h4d == _myNewVec_24_T_3[6:0] ? myVec_77 : _GEN_13430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13432 = 7'h4e == _myNewVec_24_T_3[6:0] ? myVec_78 : _GEN_13431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13433 = 7'h4f == _myNewVec_24_T_3[6:0] ? myVec_79 : _GEN_13432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13434 = 7'h50 == _myNewVec_24_T_3[6:0] ? myVec_80 : _GEN_13433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13435 = 7'h51 == _myNewVec_24_T_3[6:0] ? myVec_81 : _GEN_13434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13436 = 7'h52 == _myNewVec_24_T_3[6:0] ? myVec_82 : _GEN_13435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13437 = 7'h53 == _myNewVec_24_T_3[6:0] ? myVec_83 : _GEN_13436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13438 = 7'h54 == _myNewVec_24_T_3[6:0] ? myVec_84 : _GEN_13437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13439 = 7'h55 == _myNewVec_24_T_3[6:0] ? myVec_85 : _GEN_13438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13440 = 7'h56 == _myNewVec_24_T_3[6:0] ? myVec_86 : _GEN_13439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13441 = 7'h57 == _myNewVec_24_T_3[6:0] ? myVec_87 : _GEN_13440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13442 = 7'h58 == _myNewVec_24_T_3[6:0] ? myVec_88 : _GEN_13441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13443 = 7'h59 == _myNewVec_24_T_3[6:0] ? myVec_89 : _GEN_13442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13444 = 7'h5a == _myNewVec_24_T_3[6:0] ? myVec_90 : _GEN_13443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13445 = 7'h5b == _myNewVec_24_T_3[6:0] ? myVec_91 : _GEN_13444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13446 = 7'h5c == _myNewVec_24_T_3[6:0] ? myVec_92 : _GEN_13445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13447 = 7'h5d == _myNewVec_24_T_3[6:0] ? myVec_93 : _GEN_13446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13448 = 7'h5e == _myNewVec_24_T_3[6:0] ? myVec_94 : _GEN_13447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13449 = 7'h5f == _myNewVec_24_T_3[6:0] ? myVec_95 : _GEN_13448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13450 = 7'h60 == _myNewVec_24_T_3[6:0] ? myVec_96 : _GEN_13449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13451 = 7'h61 == _myNewVec_24_T_3[6:0] ? myVec_97 : _GEN_13450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13452 = 7'h62 == _myNewVec_24_T_3[6:0] ? myVec_98 : _GEN_13451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13453 = 7'h63 == _myNewVec_24_T_3[6:0] ? myVec_99 : _GEN_13452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13454 = 7'h64 == _myNewVec_24_T_3[6:0] ? myVec_100 : _GEN_13453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13455 = 7'h65 == _myNewVec_24_T_3[6:0] ? myVec_101 : _GEN_13454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13456 = 7'h66 == _myNewVec_24_T_3[6:0] ? myVec_102 : _GEN_13455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13457 = 7'h67 == _myNewVec_24_T_3[6:0] ? myVec_103 : _GEN_13456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13458 = 7'h68 == _myNewVec_24_T_3[6:0] ? myVec_104 : _GEN_13457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13459 = 7'h69 == _myNewVec_24_T_3[6:0] ? myVec_105 : _GEN_13458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13460 = 7'h6a == _myNewVec_24_T_3[6:0] ? myVec_106 : _GEN_13459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13461 = 7'h6b == _myNewVec_24_T_3[6:0] ? myVec_107 : _GEN_13460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13462 = 7'h6c == _myNewVec_24_T_3[6:0] ? myVec_108 : _GEN_13461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13463 = 7'h6d == _myNewVec_24_T_3[6:0] ? myVec_109 : _GEN_13462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13464 = 7'h6e == _myNewVec_24_T_3[6:0] ? myVec_110 : _GEN_13463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13465 = 7'h6f == _myNewVec_24_T_3[6:0] ? myVec_111 : _GEN_13464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13466 = 7'h70 == _myNewVec_24_T_3[6:0] ? myVec_112 : _GEN_13465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13467 = 7'h71 == _myNewVec_24_T_3[6:0] ? myVec_113 : _GEN_13466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13468 = 7'h72 == _myNewVec_24_T_3[6:0] ? myVec_114 : _GEN_13467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13469 = 7'h73 == _myNewVec_24_T_3[6:0] ? myVec_115 : _GEN_13468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13470 = 7'h74 == _myNewVec_24_T_3[6:0] ? myVec_116 : _GEN_13469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13471 = 7'h75 == _myNewVec_24_T_3[6:0] ? myVec_117 : _GEN_13470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13472 = 7'h76 == _myNewVec_24_T_3[6:0] ? myVec_118 : _GEN_13471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13473 = 7'h77 == _myNewVec_24_T_3[6:0] ? myVec_119 : _GEN_13472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13474 = 7'h78 == _myNewVec_24_T_3[6:0] ? myVec_120 : _GEN_13473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13475 = 7'h79 == _myNewVec_24_T_3[6:0] ? myVec_121 : _GEN_13474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13476 = 7'h7a == _myNewVec_24_T_3[6:0] ? myVec_122 : _GEN_13475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13477 = 7'h7b == _myNewVec_24_T_3[6:0] ? myVec_123 : _GEN_13476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13478 = 7'h7c == _myNewVec_24_T_3[6:0] ? myVec_124 : _GEN_13477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13479 = 7'h7d == _myNewVec_24_T_3[6:0] ? myVec_125 : _GEN_13478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13480 = 7'h7e == _myNewVec_24_T_3[6:0] ? myVec_126 : _GEN_13479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_24 = 7'h7f == _myNewVec_24_T_3[6:0] ? myVec_127 : _GEN_13480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_23_T_3 = _myNewVec_127_T_1 + 16'h68; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_13483 = 7'h1 == _myNewVec_23_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13484 = 7'h2 == _myNewVec_23_T_3[6:0] ? myVec_2 : _GEN_13483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13485 = 7'h3 == _myNewVec_23_T_3[6:0] ? myVec_3 : _GEN_13484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13486 = 7'h4 == _myNewVec_23_T_3[6:0] ? myVec_4 : _GEN_13485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13487 = 7'h5 == _myNewVec_23_T_3[6:0] ? myVec_5 : _GEN_13486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13488 = 7'h6 == _myNewVec_23_T_3[6:0] ? myVec_6 : _GEN_13487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13489 = 7'h7 == _myNewVec_23_T_3[6:0] ? myVec_7 : _GEN_13488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13490 = 7'h8 == _myNewVec_23_T_3[6:0] ? myVec_8 : _GEN_13489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13491 = 7'h9 == _myNewVec_23_T_3[6:0] ? myVec_9 : _GEN_13490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13492 = 7'ha == _myNewVec_23_T_3[6:0] ? myVec_10 : _GEN_13491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13493 = 7'hb == _myNewVec_23_T_3[6:0] ? myVec_11 : _GEN_13492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13494 = 7'hc == _myNewVec_23_T_3[6:0] ? myVec_12 : _GEN_13493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13495 = 7'hd == _myNewVec_23_T_3[6:0] ? myVec_13 : _GEN_13494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13496 = 7'he == _myNewVec_23_T_3[6:0] ? myVec_14 : _GEN_13495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13497 = 7'hf == _myNewVec_23_T_3[6:0] ? myVec_15 : _GEN_13496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13498 = 7'h10 == _myNewVec_23_T_3[6:0] ? myVec_16 : _GEN_13497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13499 = 7'h11 == _myNewVec_23_T_3[6:0] ? myVec_17 : _GEN_13498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13500 = 7'h12 == _myNewVec_23_T_3[6:0] ? myVec_18 : _GEN_13499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13501 = 7'h13 == _myNewVec_23_T_3[6:0] ? myVec_19 : _GEN_13500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13502 = 7'h14 == _myNewVec_23_T_3[6:0] ? myVec_20 : _GEN_13501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13503 = 7'h15 == _myNewVec_23_T_3[6:0] ? myVec_21 : _GEN_13502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13504 = 7'h16 == _myNewVec_23_T_3[6:0] ? myVec_22 : _GEN_13503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13505 = 7'h17 == _myNewVec_23_T_3[6:0] ? myVec_23 : _GEN_13504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13506 = 7'h18 == _myNewVec_23_T_3[6:0] ? myVec_24 : _GEN_13505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13507 = 7'h19 == _myNewVec_23_T_3[6:0] ? myVec_25 : _GEN_13506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13508 = 7'h1a == _myNewVec_23_T_3[6:0] ? myVec_26 : _GEN_13507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13509 = 7'h1b == _myNewVec_23_T_3[6:0] ? myVec_27 : _GEN_13508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13510 = 7'h1c == _myNewVec_23_T_3[6:0] ? myVec_28 : _GEN_13509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13511 = 7'h1d == _myNewVec_23_T_3[6:0] ? myVec_29 : _GEN_13510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13512 = 7'h1e == _myNewVec_23_T_3[6:0] ? myVec_30 : _GEN_13511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13513 = 7'h1f == _myNewVec_23_T_3[6:0] ? myVec_31 : _GEN_13512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13514 = 7'h20 == _myNewVec_23_T_3[6:0] ? myVec_32 : _GEN_13513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13515 = 7'h21 == _myNewVec_23_T_3[6:0] ? myVec_33 : _GEN_13514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13516 = 7'h22 == _myNewVec_23_T_3[6:0] ? myVec_34 : _GEN_13515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13517 = 7'h23 == _myNewVec_23_T_3[6:0] ? myVec_35 : _GEN_13516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13518 = 7'h24 == _myNewVec_23_T_3[6:0] ? myVec_36 : _GEN_13517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13519 = 7'h25 == _myNewVec_23_T_3[6:0] ? myVec_37 : _GEN_13518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13520 = 7'h26 == _myNewVec_23_T_3[6:0] ? myVec_38 : _GEN_13519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13521 = 7'h27 == _myNewVec_23_T_3[6:0] ? myVec_39 : _GEN_13520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13522 = 7'h28 == _myNewVec_23_T_3[6:0] ? myVec_40 : _GEN_13521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13523 = 7'h29 == _myNewVec_23_T_3[6:0] ? myVec_41 : _GEN_13522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13524 = 7'h2a == _myNewVec_23_T_3[6:0] ? myVec_42 : _GEN_13523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13525 = 7'h2b == _myNewVec_23_T_3[6:0] ? myVec_43 : _GEN_13524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13526 = 7'h2c == _myNewVec_23_T_3[6:0] ? myVec_44 : _GEN_13525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13527 = 7'h2d == _myNewVec_23_T_3[6:0] ? myVec_45 : _GEN_13526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13528 = 7'h2e == _myNewVec_23_T_3[6:0] ? myVec_46 : _GEN_13527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13529 = 7'h2f == _myNewVec_23_T_3[6:0] ? myVec_47 : _GEN_13528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13530 = 7'h30 == _myNewVec_23_T_3[6:0] ? myVec_48 : _GEN_13529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13531 = 7'h31 == _myNewVec_23_T_3[6:0] ? myVec_49 : _GEN_13530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13532 = 7'h32 == _myNewVec_23_T_3[6:0] ? myVec_50 : _GEN_13531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13533 = 7'h33 == _myNewVec_23_T_3[6:0] ? myVec_51 : _GEN_13532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13534 = 7'h34 == _myNewVec_23_T_3[6:0] ? myVec_52 : _GEN_13533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13535 = 7'h35 == _myNewVec_23_T_3[6:0] ? myVec_53 : _GEN_13534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13536 = 7'h36 == _myNewVec_23_T_3[6:0] ? myVec_54 : _GEN_13535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13537 = 7'h37 == _myNewVec_23_T_3[6:0] ? myVec_55 : _GEN_13536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13538 = 7'h38 == _myNewVec_23_T_3[6:0] ? myVec_56 : _GEN_13537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13539 = 7'h39 == _myNewVec_23_T_3[6:0] ? myVec_57 : _GEN_13538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13540 = 7'h3a == _myNewVec_23_T_3[6:0] ? myVec_58 : _GEN_13539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13541 = 7'h3b == _myNewVec_23_T_3[6:0] ? myVec_59 : _GEN_13540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13542 = 7'h3c == _myNewVec_23_T_3[6:0] ? myVec_60 : _GEN_13541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13543 = 7'h3d == _myNewVec_23_T_3[6:0] ? myVec_61 : _GEN_13542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13544 = 7'h3e == _myNewVec_23_T_3[6:0] ? myVec_62 : _GEN_13543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13545 = 7'h3f == _myNewVec_23_T_3[6:0] ? myVec_63 : _GEN_13544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13546 = 7'h40 == _myNewVec_23_T_3[6:0] ? myVec_64 : _GEN_13545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13547 = 7'h41 == _myNewVec_23_T_3[6:0] ? myVec_65 : _GEN_13546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13548 = 7'h42 == _myNewVec_23_T_3[6:0] ? myVec_66 : _GEN_13547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13549 = 7'h43 == _myNewVec_23_T_3[6:0] ? myVec_67 : _GEN_13548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13550 = 7'h44 == _myNewVec_23_T_3[6:0] ? myVec_68 : _GEN_13549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13551 = 7'h45 == _myNewVec_23_T_3[6:0] ? myVec_69 : _GEN_13550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13552 = 7'h46 == _myNewVec_23_T_3[6:0] ? myVec_70 : _GEN_13551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13553 = 7'h47 == _myNewVec_23_T_3[6:0] ? myVec_71 : _GEN_13552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13554 = 7'h48 == _myNewVec_23_T_3[6:0] ? myVec_72 : _GEN_13553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13555 = 7'h49 == _myNewVec_23_T_3[6:0] ? myVec_73 : _GEN_13554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13556 = 7'h4a == _myNewVec_23_T_3[6:0] ? myVec_74 : _GEN_13555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13557 = 7'h4b == _myNewVec_23_T_3[6:0] ? myVec_75 : _GEN_13556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13558 = 7'h4c == _myNewVec_23_T_3[6:0] ? myVec_76 : _GEN_13557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13559 = 7'h4d == _myNewVec_23_T_3[6:0] ? myVec_77 : _GEN_13558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13560 = 7'h4e == _myNewVec_23_T_3[6:0] ? myVec_78 : _GEN_13559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13561 = 7'h4f == _myNewVec_23_T_3[6:0] ? myVec_79 : _GEN_13560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13562 = 7'h50 == _myNewVec_23_T_3[6:0] ? myVec_80 : _GEN_13561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13563 = 7'h51 == _myNewVec_23_T_3[6:0] ? myVec_81 : _GEN_13562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13564 = 7'h52 == _myNewVec_23_T_3[6:0] ? myVec_82 : _GEN_13563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13565 = 7'h53 == _myNewVec_23_T_3[6:0] ? myVec_83 : _GEN_13564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13566 = 7'h54 == _myNewVec_23_T_3[6:0] ? myVec_84 : _GEN_13565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13567 = 7'h55 == _myNewVec_23_T_3[6:0] ? myVec_85 : _GEN_13566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13568 = 7'h56 == _myNewVec_23_T_3[6:0] ? myVec_86 : _GEN_13567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13569 = 7'h57 == _myNewVec_23_T_3[6:0] ? myVec_87 : _GEN_13568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13570 = 7'h58 == _myNewVec_23_T_3[6:0] ? myVec_88 : _GEN_13569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13571 = 7'h59 == _myNewVec_23_T_3[6:0] ? myVec_89 : _GEN_13570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13572 = 7'h5a == _myNewVec_23_T_3[6:0] ? myVec_90 : _GEN_13571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13573 = 7'h5b == _myNewVec_23_T_3[6:0] ? myVec_91 : _GEN_13572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13574 = 7'h5c == _myNewVec_23_T_3[6:0] ? myVec_92 : _GEN_13573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13575 = 7'h5d == _myNewVec_23_T_3[6:0] ? myVec_93 : _GEN_13574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13576 = 7'h5e == _myNewVec_23_T_3[6:0] ? myVec_94 : _GEN_13575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13577 = 7'h5f == _myNewVec_23_T_3[6:0] ? myVec_95 : _GEN_13576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13578 = 7'h60 == _myNewVec_23_T_3[6:0] ? myVec_96 : _GEN_13577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13579 = 7'h61 == _myNewVec_23_T_3[6:0] ? myVec_97 : _GEN_13578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13580 = 7'h62 == _myNewVec_23_T_3[6:0] ? myVec_98 : _GEN_13579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13581 = 7'h63 == _myNewVec_23_T_3[6:0] ? myVec_99 : _GEN_13580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13582 = 7'h64 == _myNewVec_23_T_3[6:0] ? myVec_100 : _GEN_13581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13583 = 7'h65 == _myNewVec_23_T_3[6:0] ? myVec_101 : _GEN_13582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13584 = 7'h66 == _myNewVec_23_T_3[6:0] ? myVec_102 : _GEN_13583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13585 = 7'h67 == _myNewVec_23_T_3[6:0] ? myVec_103 : _GEN_13584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13586 = 7'h68 == _myNewVec_23_T_3[6:0] ? myVec_104 : _GEN_13585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13587 = 7'h69 == _myNewVec_23_T_3[6:0] ? myVec_105 : _GEN_13586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13588 = 7'h6a == _myNewVec_23_T_3[6:0] ? myVec_106 : _GEN_13587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13589 = 7'h6b == _myNewVec_23_T_3[6:0] ? myVec_107 : _GEN_13588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13590 = 7'h6c == _myNewVec_23_T_3[6:0] ? myVec_108 : _GEN_13589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13591 = 7'h6d == _myNewVec_23_T_3[6:0] ? myVec_109 : _GEN_13590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13592 = 7'h6e == _myNewVec_23_T_3[6:0] ? myVec_110 : _GEN_13591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13593 = 7'h6f == _myNewVec_23_T_3[6:0] ? myVec_111 : _GEN_13592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13594 = 7'h70 == _myNewVec_23_T_3[6:0] ? myVec_112 : _GEN_13593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13595 = 7'h71 == _myNewVec_23_T_3[6:0] ? myVec_113 : _GEN_13594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13596 = 7'h72 == _myNewVec_23_T_3[6:0] ? myVec_114 : _GEN_13595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13597 = 7'h73 == _myNewVec_23_T_3[6:0] ? myVec_115 : _GEN_13596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13598 = 7'h74 == _myNewVec_23_T_3[6:0] ? myVec_116 : _GEN_13597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13599 = 7'h75 == _myNewVec_23_T_3[6:0] ? myVec_117 : _GEN_13598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13600 = 7'h76 == _myNewVec_23_T_3[6:0] ? myVec_118 : _GEN_13599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13601 = 7'h77 == _myNewVec_23_T_3[6:0] ? myVec_119 : _GEN_13600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13602 = 7'h78 == _myNewVec_23_T_3[6:0] ? myVec_120 : _GEN_13601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13603 = 7'h79 == _myNewVec_23_T_3[6:0] ? myVec_121 : _GEN_13602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13604 = 7'h7a == _myNewVec_23_T_3[6:0] ? myVec_122 : _GEN_13603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13605 = 7'h7b == _myNewVec_23_T_3[6:0] ? myVec_123 : _GEN_13604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13606 = 7'h7c == _myNewVec_23_T_3[6:0] ? myVec_124 : _GEN_13605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13607 = 7'h7d == _myNewVec_23_T_3[6:0] ? myVec_125 : _GEN_13606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13608 = 7'h7e == _myNewVec_23_T_3[6:0] ? myVec_126 : _GEN_13607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_23 = 7'h7f == _myNewVec_23_T_3[6:0] ? myVec_127 : _GEN_13608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_22_T_3 = _myNewVec_127_T_1 + 16'h69; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_13611 = 7'h1 == _myNewVec_22_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13612 = 7'h2 == _myNewVec_22_T_3[6:0] ? myVec_2 : _GEN_13611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13613 = 7'h3 == _myNewVec_22_T_3[6:0] ? myVec_3 : _GEN_13612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13614 = 7'h4 == _myNewVec_22_T_3[6:0] ? myVec_4 : _GEN_13613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13615 = 7'h5 == _myNewVec_22_T_3[6:0] ? myVec_5 : _GEN_13614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13616 = 7'h6 == _myNewVec_22_T_3[6:0] ? myVec_6 : _GEN_13615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13617 = 7'h7 == _myNewVec_22_T_3[6:0] ? myVec_7 : _GEN_13616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13618 = 7'h8 == _myNewVec_22_T_3[6:0] ? myVec_8 : _GEN_13617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13619 = 7'h9 == _myNewVec_22_T_3[6:0] ? myVec_9 : _GEN_13618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13620 = 7'ha == _myNewVec_22_T_3[6:0] ? myVec_10 : _GEN_13619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13621 = 7'hb == _myNewVec_22_T_3[6:0] ? myVec_11 : _GEN_13620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13622 = 7'hc == _myNewVec_22_T_3[6:0] ? myVec_12 : _GEN_13621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13623 = 7'hd == _myNewVec_22_T_3[6:0] ? myVec_13 : _GEN_13622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13624 = 7'he == _myNewVec_22_T_3[6:0] ? myVec_14 : _GEN_13623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13625 = 7'hf == _myNewVec_22_T_3[6:0] ? myVec_15 : _GEN_13624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13626 = 7'h10 == _myNewVec_22_T_3[6:0] ? myVec_16 : _GEN_13625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13627 = 7'h11 == _myNewVec_22_T_3[6:0] ? myVec_17 : _GEN_13626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13628 = 7'h12 == _myNewVec_22_T_3[6:0] ? myVec_18 : _GEN_13627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13629 = 7'h13 == _myNewVec_22_T_3[6:0] ? myVec_19 : _GEN_13628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13630 = 7'h14 == _myNewVec_22_T_3[6:0] ? myVec_20 : _GEN_13629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13631 = 7'h15 == _myNewVec_22_T_3[6:0] ? myVec_21 : _GEN_13630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13632 = 7'h16 == _myNewVec_22_T_3[6:0] ? myVec_22 : _GEN_13631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13633 = 7'h17 == _myNewVec_22_T_3[6:0] ? myVec_23 : _GEN_13632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13634 = 7'h18 == _myNewVec_22_T_3[6:0] ? myVec_24 : _GEN_13633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13635 = 7'h19 == _myNewVec_22_T_3[6:0] ? myVec_25 : _GEN_13634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13636 = 7'h1a == _myNewVec_22_T_3[6:0] ? myVec_26 : _GEN_13635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13637 = 7'h1b == _myNewVec_22_T_3[6:0] ? myVec_27 : _GEN_13636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13638 = 7'h1c == _myNewVec_22_T_3[6:0] ? myVec_28 : _GEN_13637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13639 = 7'h1d == _myNewVec_22_T_3[6:0] ? myVec_29 : _GEN_13638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13640 = 7'h1e == _myNewVec_22_T_3[6:0] ? myVec_30 : _GEN_13639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13641 = 7'h1f == _myNewVec_22_T_3[6:0] ? myVec_31 : _GEN_13640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13642 = 7'h20 == _myNewVec_22_T_3[6:0] ? myVec_32 : _GEN_13641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13643 = 7'h21 == _myNewVec_22_T_3[6:0] ? myVec_33 : _GEN_13642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13644 = 7'h22 == _myNewVec_22_T_3[6:0] ? myVec_34 : _GEN_13643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13645 = 7'h23 == _myNewVec_22_T_3[6:0] ? myVec_35 : _GEN_13644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13646 = 7'h24 == _myNewVec_22_T_3[6:0] ? myVec_36 : _GEN_13645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13647 = 7'h25 == _myNewVec_22_T_3[6:0] ? myVec_37 : _GEN_13646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13648 = 7'h26 == _myNewVec_22_T_3[6:0] ? myVec_38 : _GEN_13647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13649 = 7'h27 == _myNewVec_22_T_3[6:0] ? myVec_39 : _GEN_13648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13650 = 7'h28 == _myNewVec_22_T_3[6:0] ? myVec_40 : _GEN_13649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13651 = 7'h29 == _myNewVec_22_T_3[6:0] ? myVec_41 : _GEN_13650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13652 = 7'h2a == _myNewVec_22_T_3[6:0] ? myVec_42 : _GEN_13651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13653 = 7'h2b == _myNewVec_22_T_3[6:0] ? myVec_43 : _GEN_13652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13654 = 7'h2c == _myNewVec_22_T_3[6:0] ? myVec_44 : _GEN_13653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13655 = 7'h2d == _myNewVec_22_T_3[6:0] ? myVec_45 : _GEN_13654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13656 = 7'h2e == _myNewVec_22_T_3[6:0] ? myVec_46 : _GEN_13655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13657 = 7'h2f == _myNewVec_22_T_3[6:0] ? myVec_47 : _GEN_13656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13658 = 7'h30 == _myNewVec_22_T_3[6:0] ? myVec_48 : _GEN_13657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13659 = 7'h31 == _myNewVec_22_T_3[6:0] ? myVec_49 : _GEN_13658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13660 = 7'h32 == _myNewVec_22_T_3[6:0] ? myVec_50 : _GEN_13659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13661 = 7'h33 == _myNewVec_22_T_3[6:0] ? myVec_51 : _GEN_13660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13662 = 7'h34 == _myNewVec_22_T_3[6:0] ? myVec_52 : _GEN_13661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13663 = 7'h35 == _myNewVec_22_T_3[6:0] ? myVec_53 : _GEN_13662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13664 = 7'h36 == _myNewVec_22_T_3[6:0] ? myVec_54 : _GEN_13663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13665 = 7'h37 == _myNewVec_22_T_3[6:0] ? myVec_55 : _GEN_13664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13666 = 7'h38 == _myNewVec_22_T_3[6:0] ? myVec_56 : _GEN_13665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13667 = 7'h39 == _myNewVec_22_T_3[6:0] ? myVec_57 : _GEN_13666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13668 = 7'h3a == _myNewVec_22_T_3[6:0] ? myVec_58 : _GEN_13667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13669 = 7'h3b == _myNewVec_22_T_3[6:0] ? myVec_59 : _GEN_13668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13670 = 7'h3c == _myNewVec_22_T_3[6:0] ? myVec_60 : _GEN_13669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13671 = 7'h3d == _myNewVec_22_T_3[6:0] ? myVec_61 : _GEN_13670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13672 = 7'h3e == _myNewVec_22_T_3[6:0] ? myVec_62 : _GEN_13671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13673 = 7'h3f == _myNewVec_22_T_3[6:0] ? myVec_63 : _GEN_13672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13674 = 7'h40 == _myNewVec_22_T_3[6:0] ? myVec_64 : _GEN_13673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13675 = 7'h41 == _myNewVec_22_T_3[6:0] ? myVec_65 : _GEN_13674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13676 = 7'h42 == _myNewVec_22_T_3[6:0] ? myVec_66 : _GEN_13675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13677 = 7'h43 == _myNewVec_22_T_3[6:0] ? myVec_67 : _GEN_13676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13678 = 7'h44 == _myNewVec_22_T_3[6:0] ? myVec_68 : _GEN_13677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13679 = 7'h45 == _myNewVec_22_T_3[6:0] ? myVec_69 : _GEN_13678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13680 = 7'h46 == _myNewVec_22_T_3[6:0] ? myVec_70 : _GEN_13679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13681 = 7'h47 == _myNewVec_22_T_3[6:0] ? myVec_71 : _GEN_13680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13682 = 7'h48 == _myNewVec_22_T_3[6:0] ? myVec_72 : _GEN_13681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13683 = 7'h49 == _myNewVec_22_T_3[6:0] ? myVec_73 : _GEN_13682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13684 = 7'h4a == _myNewVec_22_T_3[6:0] ? myVec_74 : _GEN_13683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13685 = 7'h4b == _myNewVec_22_T_3[6:0] ? myVec_75 : _GEN_13684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13686 = 7'h4c == _myNewVec_22_T_3[6:0] ? myVec_76 : _GEN_13685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13687 = 7'h4d == _myNewVec_22_T_3[6:0] ? myVec_77 : _GEN_13686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13688 = 7'h4e == _myNewVec_22_T_3[6:0] ? myVec_78 : _GEN_13687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13689 = 7'h4f == _myNewVec_22_T_3[6:0] ? myVec_79 : _GEN_13688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13690 = 7'h50 == _myNewVec_22_T_3[6:0] ? myVec_80 : _GEN_13689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13691 = 7'h51 == _myNewVec_22_T_3[6:0] ? myVec_81 : _GEN_13690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13692 = 7'h52 == _myNewVec_22_T_3[6:0] ? myVec_82 : _GEN_13691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13693 = 7'h53 == _myNewVec_22_T_3[6:0] ? myVec_83 : _GEN_13692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13694 = 7'h54 == _myNewVec_22_T_3[6:0] ? myVec_84 : _GEN_13693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13695 = 7'h55 == _myNewVec_22_T_3[6:0] ? myVec_85 : _GEN_13694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13696 = 7'h56 == _myNewVec_22_T_3[6:0] ? myVec_86 : _GEN_13695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13697 = 7'h57 == _myNewVec_22_T_3[6:0] ? myVec_87 : _GEN_13696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13698 = 7'h58 == _myNewVec_22_T_3[6:0] ? myVec_88 : _GEN_13697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13699 = 7'h59 == _myNewVec_22_T_3[6:0] ? myVec_89 : _GEN_13698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13700 = 7'h5a == _myNewVec_22_T_3[6:0] ? myVec_90 : _GEN_13699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13701 = 7'h5b == _myNewVec_22_T_3[6:0] ? myVec_91 : _GEN_13700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13702 = 7'h5c == _myNewVec_22_T_3[6:0] ? myVec_92 : _GEN_13701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13703 = 7'h5d == _myNewVec_22_T_3[6:0] ? myVec_93 : _GEN_13702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13704 = 7'h5e == _myNewVec_22_T_3[6:0] ? myVec_94 : _GEN_13703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13705 = 7'h5f == _myNewVec_22_T_3[6:0] ? myVec_95 : _GEN_13704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13706 = 7'h60 == _myNewVec_22_T_3[6:0] ? myVec_96 : _GEN_13705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13707 = 7'h61 == _myNewVec_22_T_3[6:0] ? myVec_97 : _GEN_13706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13708 = 7'h62 == _myNewVec_22_T_3[6:0] ? myVec_98 : _GEN_13707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13709 = 7'h63 == _myNewVec_22_T_3[6:0] ? myVec_99 : _GEN_13708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13710 = 7'h64 == _myNewVec_22_T_3[6:0] ? myVec_100 : _GEN_13709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13711 = 7'h65 == _myNewVec_22_T_3[6:0] ? myVec_101 : _GEN_13710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13712 = 7'h66 == _myNewVec_22_T_3[6:0] ? myVec_102 : _GEN_13711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13713 = 7'h67 == _myNewVec_22_T_3[6:0] ? myVec_103 : _GEN_13712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13714 = 7'h68 == _myNewVec_22_T_3[6:0] ? myVec_104 : _GEN_13713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13715 = 7'h69 == _myNewVec_22_T_3[6:0] ? myVec_105 : _GEN_13714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13716 = 7'h6a == _myNewVec_22_T_3[6:0] ? myVec_106 : _GEN_13715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13717 = 7'h6b == _myNewVec_22_T_3[6:0] ? myVec_107 : _GEN_13716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13718 = 7'h6c == _myNewVec_22_T_3[6:0] ? myVec_108 : _GEN_13717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13719 = 7'h6d == _myNewVec_22_T_3[6:0] ? myVec_109 : _GEN_13718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13720 = 7'h6e == _myNewVec_22_T_3[6:0] ? myVec_110 : _GEN_13719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13721 = 7'h6f == _myNewVec_22_T_3[6:0] ? myVec_111 : _GEN_13720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13722 = 7'h70 == _myNewVec_22_T_3[6:0] ? myVec_112 : _GEN_13721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13723 = 7'h71 == _myNewVec_22_T_3[6:0] ? myVec_113 : _GEN_13722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13724 = 7'h72 == _myNewVec_22_T_3[6:0] ? myVec_114 : _GEN_13723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13725 = 7'h73 == _myNewVec_22_T_3[6:0] ? myVec_115 : _GEN_13724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13726 = 7'h74 == _myNewVec_22_T_3[6:0] ? myVec_116 : _GEN_13725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13727 = 7'h75 == _myNewVec_22_T_3[6:0] ? myVec_117 : _GEN_13726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13728 = 7'h76 == _myNewVec_22_T_3[6:0] ? myVec_118 : _GEN_13727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13729 = 7'h77 == _myNewVec_22_T_3[6:0] ? myVec_119 : _GEN_13728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13730 = 7'h78 == _myNewVec_22_T_3[6:0] ? myVec_120 : _GEN_13729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13731 = 7'h79 == _myNewVec_22_T_3[6:0] ? myVec_121 : _GEN_13730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13732 = 7'h7a == _myNewVec_22_T_3[6:0] ? myVec_122 : _GEN_13731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13733 = 7'h7b == _myNewVec_22_T_3[6:0] ? myVec_123 : _GEN_13732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13734 = 7'h7c == _myNewVec_22_T_3[6:0] ? myVec_124 : _GEN_13733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13735 = 7'h7d == _myNewVec_22_T_3[6:0] ? myVec_125 : _GEN_13734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13736 = 7'h7e == _myNewVec_22_T_3[6:0] ? myVec_126 : _GEN_13735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_22 = 7'h7f == _myNewVec_22_T_3[6:0] ? myVec_127 : _GEN_13736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_21_T_3 = _myNewVec_127_T_1 + 16'h6a; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_13739 = 7'h1 == _myNewVec_21_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13740 = 7'h2 == _myNewVec_21_T_3[6:0] ? myVec_2 : _GEN_13739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13741 = 7'h3 == _myNewVec_21_T_3[6:0] ? myVec_3 : _GEN_13740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13742 = 7'h4 == _myNewVec_21_T_3[6:0] ? myVec_4 : _GEN_13741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13743 = 7'h5 == _myNewVec_21_T_3[6:0] ? myVec_5 : _GEN_13742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13744 = 7'h6 == _myNewVec_21_T_3[6:0] ? myVec_6 : _GEN_13743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13745 = 7'h7 == _myNewVec_21_T_3[6:0] ? myVec_7 : _GEN_13744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13746 = 7'h8 == _myNewVec_21_T_3[6:0] ? myVec_8 : _GEN_13745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13747 = 7'h9 == _myNewVec_21_T_3[6:0] ? myVec_9 : _GEN_13746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13748 = 7'ha == _myNewVec_21_T_3[6:0] ? myVec_10 : _GEN_13747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13749 = 7'hb == _myNewVec_21_T_3[6:0] ? myVec_11 : _GEN_13748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13750 = 7'hc == _myNewVec_21_T_3[6:0] ? myVec_12 : _GEN_13749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13751 = 7'hd == _myNewVec_21_T_3[6:0] ? myVec_13 : _GEN_13750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13752 = 7'he == _myNewVec_21_T_3[6:0] ? myVec_14 : _GEN_13751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13753 = 7'hf == _myNewVec_21_T_3[6:0] ? myVec_15 : _GEN_13752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13754 = 7'h10 == _myNewVec_21_T_3[6:0] ? myVec_16 : _GEN_13753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13755 = 7'h11 == _myNewVec_21_T_3[6:0] ? myVec_17 : _GEN_13754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13756 = 7'h12 == _myNewVec_21_T_3[6:0] ? myVec_18 : _GEN_13755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13757 = 7'h13 == _myNewVec_21_T_3[6:0] ? myVec_19 : _GEN_13756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13758 = 7'h14 == _myNewVec_21_T_3[6:0] ? myVec_20 : _GEN_13757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13759 = 7'h15 == _myNewVec_21_T_3[6:0] ? myVec_21 : _GEN_13758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13760 = 7'h16 == _myNewVec_21_T_3[6:0] ? myVec_22 : _GEN_13759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13761 = 7'h17 == _myNewVec_21_T_3[6:0] ? myVec_23 : _GEN_13760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13762 = 7'h18 == _myNewVec_21_T_3[6:0] ? myVec_24 : _GEN_13761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13763 = 7'h19 == _myNewVec_21_T_3[6:0] ? myVec_25 : _GEN_13762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13764 = 7'h1a == _myNewVec_21_T_3[6:0] ? myVec_26 : _GEN_13763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13765 = 7'h1b == _myNewVec_21_T_3[6:0] ? myVec_27 : _GEN_13764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13766 = 7'h1c == _myNewVec_21_T_3[6:0] ? myVec_28 : _GEN_13765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13767 = 7'h1d == _myNewVec_21_T_3[6:0] ? myVec_29 : _GEN_13766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13768 = 7'h1e == _myNewVec_21_T_3[6:0] ? myVec_30 : _GEN_13767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13769 = 7'h1f == _myNewVec_21_T_3[6:0] ? myVec_31 : _GEN_13768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13770 = 7'h20 == _myNewVec_21_T_3[6:0] ? myVec_32 : _GEN_13769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13771 = 7'h21 == _myNewVec_21_T_3[6:0] ? myVec_33 : _GEN_13770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13772 = 7'h22 == _myNewVec_21_T_3[6:0] ? myVec_34 : _GEN_13771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13773 = 7'h23 == _myNewVec_21_T_3[6:0] ? myVec_35 : _GEN_13772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13774 = 7'h24 == _myNewVec_21_T_3[6:0] ? myVec_36 : _GEN_13773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13775 = 7'h25 == _myNewVec_21_T_3[6:0] ? myVec_37 : _GEN_13774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13776 = 7'h26 == _myNewVec_21_T_3[6:0] ? myVec_38 : _GEN_13775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13777 = 7'h27 == _myNewVec_21_T_3[6:0] ? myVec_39 : _GEN_13776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13778 = 7'h28 == _myNewVec_21_T_3[6:0] ? myVec_40 : _GEN_13777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13779 = 7'h29 == _myNewVec_21_T_3[6:0] ? myVec_41 : _GEN_13778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13780 = 7'h2a == _myNewVec_21_T_3[6:0] ? myVec_42 : _GEN_13779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13781 = 7'h2b == _myNewVec_21_T_3[6:0] ? myVec_43 : _GEN_13780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13782 = 7'h2c == _myNewVec_21_T_3[6:0] ? myVec_44 : _GEN_13781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13783 = 7'h2d == _myNewVec_21_T_3[6:0] ? myVec_45 : _GEN_13782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13784 = 7'h2e == _myNewVec_21_T_3[6:0] ? myVec_46 : _GEN_13783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13785 = 7'h2f == _myNewVec_21_T_3[6:0] ? myVec_47 : _GEN_13784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13786 = 7'h30 == _myNewVec_21_T_3[6:0] ? myVec_48 : _GEN_13785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13787 = 7'h31 == _myNewVec_21_T_3[6:0] ? myVec_49 : _GEN_13786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13788 = 7'h32 == _myNewVec_21_T_3[6:0] ? myVec_50 : _GEN_13787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13789 = 7'h33 == _myNewVec_21_T_3[6:0] ? myVec_51 : _GEN_13788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13790 = 7'h34 == _myNewVec_21_T_3[6:0] ? myVec_52 : _GEN_13789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13791 = 7'h35 == _myNewVec_21_T_3[6:0] ? myVec_53 : _GEN_13790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13792 = 7'h36 == _myNewVec_21_T_3[6:0] ? myVec_54 : _GEN_13791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13793 = 7'h37 == _myNewVec_21_T_3[6:0] ? myVec_55 : _GEN_13792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13794 = 7'h38 == _myNewVec_21_T_3[6:0] ? myVec_56 : _GEN_13793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13795 = 7'h39 == _myNewVec_21_T_3[6:0] ? myVec_57 : _GEN_13794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13796 = 7'h3a == _myNewVec_21_T_3[6:0] ? myVec_58 : _GEN_13795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13797 = 7'h3b == _myNewVec_21_T_3[6:0] ? myVec_59 : _GEN_13796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13798 = 7'h3c == _myNewVec_21_T_3[6:0] ? myVec_60 : _GEN_13797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13799 = 7'h3d == _myNewVec_21_T_3[6:0] ? myVec_61 : _GEN_13798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13800 = 7'h3e == _myNewVec_21_T_3[6:0] ? myVec_62 : _GEN_13799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13801 = 7'h3f == _myNewVec_21_T_3[6:0] ? myVec_63 : _GEN_13800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13802 = 7'h40 == _myNewVec_21_T_3[6:0] ? myVec_64 : _GEN_13801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13803 = 7'h41 == _myNewVec_21_T_3[6:0] ? myVec_65 : _GEN_13802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13804 = 7'h42 == _myNewVec_21_T_3[6:0] ? myVec_66 : _GEN_13803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13805 = 7'h43 == _myNewVec_21_T_3[6:0] ? myVec_67 : _GEN_13804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13806 = 7'h44 == _myNewVec_21_T_3[6:0] ? myVec_68 : _GEN_13805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13807 = 7'h45 == _myNewVec_21_T_3[6:0] ? myVec_69 : _GEN_13806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13808 = 7'h46 == _myNewVec_21_T_3[6:0] ? myVec_70 : _GEN_13807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13809 = 7'h47 == _myNewVec_21_T_3[6:0] ? myVec_71 : _GEN_13808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13810 = 7'h48 == _myNewVec_21_T_3[6:0] ? myVec_72 : _GEN_13809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13811 = 7'h49 == _myNewVec_21_T_3[6:0] ? myVec_73 : _GEN_13810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13812 = 7'h4a == _myNewVec_21_T_3[6:0] ? myVec_74 : _GEN_13811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13813 = 7'h4b == _myNewVec_21_T_3[6:0] ? myVec_75 : _GEN_13812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13814 = 7'h4c == _myNewVec_21_T_3[6:0] ? myVec_76 : _GEN_13813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13815 = 7'h4d == _myNewVec_21_T_3[6:0] ? myVec_77 : _GEN_13814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13816 = 7'h4e == _myNewVec_21_T_3[6:0] ? myVec_78 : _GEN_13815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13817 = 7'h4f == _myNewVec_21_T_3[6:0] ? myVec_79 : _GEN_13816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13818 = 7'h50 == _myNewVec_21_T_3[6:0] ? myVec_80 : _GEN_13817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13819 = 7'h51 == _myNewVec_21_T_3[6:0] ? myVec_81 : _GEN_13818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13820 = 7'h52 == _myNewVec_21_T_3[6:0] ? myVec_82 : _GEN_13819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13821 = 7'h53 == _myNewVec_21_T_3[6:0] ? myVec_83 : _GEN_13820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13822 = 7'h54 == _myNewVec_21_T_3[6:0] ? myVec_84 : _GEN_13821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13823 = 7'h55 == _myNewVec_21_T_3[6:0] ? myVec_85 : _GEN_13822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13824 = 7'h56 == _myNewVec_21_T_3[6:0] ? myVec_86 : _GEN_13823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13825 = 7'h57 == _myNewVec_21_T_3[6:0] ? myVec_87 : _GEN_13824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13826 = 7'h58 == _myNewVec_21_T_3[6:0] ? myVec_88 : _GEN_13825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13827 = 7'h59 == _myNewVec_21_T_3[6:0] ? myVec_89 : _GEN_13826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13828 = 7'h5a == _myNewVec_21_T_3[6:0] ? myVec_90 : _GEN_13827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13829 = 7'h5b == _myNewVec_21_T_3[6:0] ? myVec_91 : _GEN_13828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13830 = 7'h5c == _myNewVec_21_T_3[6:0] ? myVec_92 : _GEN_13829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13831 = 7'h5d == _myNewVec_21_T_3[6:0] ? myVec_93 : _GEN_13830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13832 = 7'h5e == _myNewVec_21_T_3[6:0] ? myVec_94 : _GEN_13831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13833 = 7'h5f == _myNewVec_21_T_3[6:0] ? myVec_95 : _GEN_13832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13834 = 7'h60 == _myNewVec_21_T_3[6:0] ? myVec_96 : _GEN_13833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13835 = 7'h61 == _myNewVec_21_T_3[6:0] ? myVec_97 : _GEN_13834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13836 = 7'h62 == _myNewVec_21_T_3[6:0] ? myVec_98 : _GEN_13835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13837 = 7'h63 == _myNewVec_21_T_3[6:0] ? myVec_99 : _GEN_13836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13838 = 7'h64 == _myNewVec_21_T_3[6:0] ? myVec_100 : _GEN_13837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13839 = 7'h65 == _myNewVec_21_T_3[6:0] ? myVec_101 : _GEN_13838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13840 = 7'h66 == _myNewVec_21_T_3[6:0] ? myVec_102 : _GEN_13839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13841 = 7'h67 == _myNewVec_21_T_3[6:0] ? myVec_103 : _GEN_13840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13842 = 7'h68 == _myNewVec_21_T_3[6:0] ? myVec_104 : _GEN_13841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13843 = 7'h69 == _myNewVec_21_T_3[6:0] ? myVec_105 : _GEN_13842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13844 = 7'h6a == _myNewVec_21_T_3[6:0] ? myVec_106 : _GEN_13843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13845 = 7'h6b == _myNewVec_21_T_3[6:0] ? myVec_107 : _GEN_13844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13846 = 7'h6c == _myNewVec_21_T_3[6:0] ? myVec_108 : _GEN_13845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13847 = 7'h6d == _myNewVec_21_T_3[6:0] ? myVec_109 : _GEN_13846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13848 = 7'h6e == _myNewVec_21_T_3[6:0] ? myVec_110 : _GEN_13847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13849 = 7'h6f == _myNewVec_21_T_3[6:0] ? myVec_111 : _GEN_13848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13850 = 7'h70 == _myNewVec_21_T_3[6:0] ? myVec_112 : _GEN_13849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13851 = 7'h71 == _myNewVec_21_T_3[6:0] ? myVec_113 : _GEN_13850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13852 = 7'h72 == _myNewVec_21_T_3[6:0] ? myVec_114 : _GEN_13851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13853 = 7'h73 == _myNewVec_21_T_3[6:0] ? myVec_115 : _GEN_13852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13854 = 7'h74 == _myNewVec_21_T_3[6:0] ? myVec_116 : _GEN_13853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13855 = 7'h75 == _myNewVec_21_T_3[6:0] ? myVec_117 : _GEN_13854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13856 = 7'h76 == _myNewVec_21_T_3[6:0] ? myVec_118 : _GEN_13855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13857 = 7'h77 == _myNewVec_21_T_3[6:0] ? myVec_119 : _GEN_13856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13858 = 7'h78 == _myNewVec_21_T_3[6:0] ? myVec_120 : _GEN_13857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13859 = 7'h79 == _myNewVec_21_T_3[6:0] ? myVec_121 : _GEN_13858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13860 = 7'h7a == _myNewVec_21_T_3[6:0] ? myVec_122 : _GEN_13859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13861 = 7'h7b == _myNewVec_21_T_3[6:0] ? myVec_123 : _GEN_13860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13862 = 7'h7c == _myNewVec_21_T_3[6:0] ? myVec_124 : _GEN_13861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13863 = 7'h7d == _myNewVec_21_T_3[6:0] ? myVec_125 : _GEN_13862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13864 = 7'h7e == _myNewVec_21_T_3[6:0] ? myVec_126 : _GEN_13863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_21 = 7'h7f == _myNewVec_21_T_3[6:0] ? myVec_127 : _GEN_13864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_20_T_3 = _myNewVec_127_T_1 + 16'h6b; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_13867 = 7'h1 == _myNewVec_20_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13868 = 7'h2 == _myNewVec_20_T_3[6:0] ? myVec_2 : _GEN_13867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13869 = 7'h3 == _myNewVec_20_T_3[6:0] ? myVec_3 : _GEN_13868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13870 = 7'h4 == _myNewVec_20_T_3[6:0] ? myVec_4 : _GEN_13869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13871 = 7'h5 == _myNewVec_20_T_3[6:0] ? myVec_5 : _GEN_13870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13872 = 7'h6 == _myNewVec_20_T_3[6:0] ? myVec_6 : _GEN_13871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13873 = 7'h7 == _myNewVec_20_T_3[6:0] ? myVec_7 : _GEN_13872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13874 = 7'h8 == _myNewVec_20_T_3[6:0] ? myVec_8 : _GEN_13873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13875 = 7'h9 == _myNewVec_20_T_3[6:0] ? myVec_9 : _GEN_13874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13876 = 7'ha == _myNewVec_20_T_3[6:0] ? myVec_10 : _GEN_13875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13877 = 7'hb == _myNewVec_20_T_3[6:0] ? myVec_11 : _GEN_13876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13878 = 7'hc == _myNewVec_20_T_3[6:0] ? myVec_12 : _GEN_13877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13879 = 7'hd == _myNewVec_20_T_3[6:0] ? myVec_13 : _GEN_13878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13880 = 7'he == _myNewVec_20_T_3[6:0] ? myVec_14 : _GEN_13879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13881 = 7'hf == _myNewVec_20_T_3[6:0] ? myVec_15 : _GEN_13880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13882 = 7'h10 == _myNewVec_20_T_3[6:0] ? myVec_16 : _GEN_13881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13883 = 7'h11 == _myNewVec_20_T_3[6:0] ? myVec_17 : _GEN_13882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13884 = 7'h12 == _myNewVec_20_T_3[6:0] ? myVec_18 : _GEN_13883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13885 = 7'h13 == _myNewVec_20_T_3[6:0] ? myVec_19 : _GEN_13884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13886 = 7'h14 == _myNewVec_20_T_3[6:0] ? myVec_20 : _GEN_13885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13887 = 7'h15 == _myNewVec_20_T_3[6:0] ? myVec_21 : _GEN_13886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13888 = 7'h16 == _myNewVec_20_T_3[6:0] ? myVec_22 : _GEN_13887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13889 = 7'h17 == _myNewVec_20_T_3[6:0] ? myVec_23 : _GEN_13888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13890 = 7'h18 == _myNewVec_20_T_3[6:0] ? myVec_24 : _GEN_13889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13891 = 7'h19 == _myNewVec_20_T_3[6:0] ? myVec_25 : _GEN_13890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13892 = 7'h1a == _myNewVec_20_T_3[6:0] ? myVec_26 : _GEN_13891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13893 = 7'h1b == _myNewVec_20_T_3[6:0] ? myVec_27 : _GEN_13892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13894 = 7'h1c == _myNewVec_20_T_3[6:0] ? myVec_28 : _GEN_13893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13895 = 7'h1d == _myNewVec_20_T_3[6:0] ? myVec_29 : _GEN_13894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13896 = 7'h1e == _myNewVec_20_T_3[6:0] ? myVec_30 : _GEN_13895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13897 = 7'h1f == _myNewVec_20_T_3[6:0] ? myVec_31 : _GEN_13896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13898 = 7'h20 == _myNewVec_20_T_3[6:0] ? myVec_32 : _GEN_13897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13899 = 7'h21 == _myNewVec_20_T_3[6:0] ? myVec_33 : _GEN_13898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13900 = 7'h22 == _myNewVec_20_T_3[6:0] ? myVec_34 : _GEN_13899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13901 = 7'h23 == _myNewVec_20_T_3[6:0] ? myVec_35 : _GEN_13900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13902 = 7'h24 == _myNewVec_20_T_3[6:0] ? myVec_36 : _GEN_13901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13903 = 7'h25 == _myNewVec_20_T_3[6:0] ? myVec_37 : _GEN_13902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13904 = 7'h26 == _myNewVec_20_T_3[6:0] ? myVec_38 : _GEN_13903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13905 = 7'h27 == _myNewVec_20_T_3[6:0] ? myVec_39 : _GEN_13904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13906 = 7'h28 == _myNewVec_20_T_3[6:0] ? myVec_40 : _GEN_13905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13907 = 7'h29 == _myNewVec_20_T_3[6:0] ? myVec_41 : _GEN_13906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13908 = 7'h2a == _myNewVec_20_T_3[6:0] ? myVec_42 : _GEN_13907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13909 = 7'h2b == _myNewVec_20_T_3[6:0] ? myVec_43 : _GEN_13908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13910 = 7'h2c == _myNewVec_20_T_3[6:0] ? myVec_44 : _GEN_13909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13911 = 7'h2d == _myNewVec_20_T_3[6:0] ? myVec_45 : _GEN_13910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13912 = 7'h2e == _myNewVec_20_T_3[6:0] ? myVec_46 : _GEN_13911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13913 = 7'h2f == _myNewVec_20_T_3[6:0] ? myVec_47 : _GEN_13912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13914 = 7'h30 == _myNewVec_20_T_3[6:0] ? myVec_48 : _GEN_13913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13915 = 7'h31 == _myNewVec_20_T_3[6:0] ? myVec_49 : _GEN_13914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13916 = 7'h32 == _myNewVec_20_T_3[6:0] ? myVec_50 : _GEN_13915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13917 = 7'h33 == _myNewVec_20_T_3[6:0] ? myVec_51 : _GEN_13916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13918 = 7'h34 == _myNewVec_20_T_3[6:0] ? myVec_52 : _GEN_13917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13919 = 7'h35 == _myNewVec_20_T_3[6:0] ? myVec_53 : _GEN_13918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13920 = 7'h36 == _myNewVec_20_T_3[6:0] ? myVec_54 : _GEN_13919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13921 = 7'h37 == _myNewVec_20_T_3[6:0] ? myVec_55 : _GEN_13920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13922 = 7'h38 == _myNewVec_20_T_3[6:0] ? myVec_56 : _GEN_13921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13923 = 7'h39 == _myNewVec_20_T_3[6:0] ? myVec_57 : _GEN_13922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13924 = 7'h3a == _myNewVec_20_T_3[6:0] ? myVec_58 : _GEN_13923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13925 = 7'h3b == _myNewVec_20_T_3[6:0] ? myVec_59 : _GEN_13924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13926 = 7'h3c == _myNewVec_20_T_3[6:0] ? myVec_60 : _GEN_13925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13927 = 7'h3d == _myNewVec_20_T_3[6:0] ? myVec_61 : _GEN_13926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13928 = 7'h3e == _myNewVec_20_T_3[6:0] ? myVec_62 : _GEN_13927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13929 = 7'h3f == _myNewVec_20_T_3[6:0] ? myVec_63 : _GEN_13928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13930 = 7'h40 == _myNewVec_20_T_3[6:0] ? myVec_64 : _GEN_13929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13931 = 7'h41 == _myNewVec_20_T_3[6:0] ? myVec_65 : _GEN_13930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13932 = 7'h42 == _myNewVec_20_T_3[6:0] ? myVec_66 : _GEN_13931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13933 = 7'h43 == _myNewVec_20_T_3[6:0] ? myVec_67 : _GEN_13932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13934 = 7'h44 == _myNewVec_20_T_3[6:0] ? myVec_68 : _GEN_13933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13935 = 7'h45 == _myNewVec_20_T_3[6:0] ? myVec_69 : _GEN_13934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13936 = 7'h46 == _myNewVec_20_T_3[6:0] ? myVec_70 : _GEN_13935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13937 = 7'h47 == _myNewVec_20_T_3[6:0] ? myVec_71 : _GEN_13936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13938 = 7'h48 == _myNewVec_20_T_3[6:0] ? myVec_72 : _GEN_13937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13939 = 7'h49 == _myNewVec_20_T_3[6:0] ? myVec_73 : _GEN_13938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13940 = 7'h4a == _myNewVec_20_T_3[6:0] ? myVec_74 : _GEN_13939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13941 = 7'h4b == _myNewVec_20_T_3[6:0] ? myVec_75 : _GEN_13940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13942 = 7'h4c == _myNewVec_20_T_3[6:0] ? myVec_76 : _GEN_13941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13943 = 7'h4d == _myNewVec_20_T_3[6:0] ? myVec_77 : _GEN_13942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13944 = 7'h4e == _myNewVec_20_T_3[6:0] ? myVec_78 : _GEN_13943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13945 = 7'h4f == _myNewVec_20_T_3[6:0] ? myVec_79 : _GEN_13944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13946 = 7'h50 == _myNewVec_20_T_3[6:0] ? myVec_80 : _GEN_13945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13947 = 7'h51 == _myNewVec_20_T_3[6:0] ? myVec_81 : _GEN_13946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13948 = 7'h52 == _myNewVec_20_T_3[6:0] ? myVec_82 : _GEN_13947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13949 = 7'h53 == _myNewVec_20_T_3[6:0] ? myVec_83 : _GEN_13948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13950 = 7'h54 == _myNewVec_20_T_3[6:0] ? myVec_84 : _GEN_13949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13951 = 7'h55 == _myNewVec_20_T_3[6:0] ? myVec_85 : _GEN_13950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13952 = 7'h56 == _myNewVec_20_T_3[6:0] ? myVec_86 : _GEN_13951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13953 = 7'h57 == _myNewVec_20_T_3[6:0] ? myVec_87 : _GEN_13952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13954 = 7'h58 == _myNewVec_20_T_3[6:0] ? myVec_88 : _GEN_13953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13955 = 7'h59 == _myNewVec_20_T_3[6:0] ? myVec_89 : _GEN_13954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13956 = 7'h5a == _myNewVec_20_T_3[6:0] ? myVec_90 : _GEN_13955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13957 = 7'h5b == _myNewVec_20_T_3[6:0] ? myVec_91 : _GEN_13956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13958 = 7'h5c == _myNewVec_20_T_3[6:0] ? myVec_92 : _GEN_13957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13959 = 7'h5d == _myNewVec_20_T_3[6:0] ? myVec_93 : _GEN_13958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13960 = 7'h5e == _myNewVec_20_T_3[6:0] ? myVec_94 : _GEN_13959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13961 = 7'h5f == _myNewVec_20_T_3[6:0] ? myVec_95 : _GEN_13960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13962 = 7'h60 == _myNewVec_20_T_3[6:0] ? myVec_96 : _GEN_13961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13963 = 7'h61 == _myNewVec_20_T_3[6:0] ? myVec_97 : _GEN_13962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13964 = 7'h62 == _myNewVec_20_T_3[6:0] ? myVec_98 : _GEN_13963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13965 = 7'h63 == _myNewVec_20_T_3[6:0] ? myVec_99 : _GEN_13964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13966 = 7'h64 == _myNewVec_20_T_3[6:0] ? myVec_100 : _GEN_13965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13967 = 7'h65 == _myNewVec_20_T_3[6:0] ? myVec_101 : _GEN_13966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13968 = 7'h66 == _myNewVec_20_T_3[6:0] ? myVec_102 : _GEN_13967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13969 = 7'h67 == _myNewVec_20_T_3[6:0] ? myVec_103 : _GEN_13968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13970 = 7'h68 == _myNewVec_20_T_3[6:0] ? myVec_104 : _GEN_13969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13971 = 7'h69 == _myNewVec_20_T_3[6:0] ? myVec_105 : _GEN_13970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13972 = 7'h6a == _myNewVec_20_T_3[6:0] ? myVec_106 : _GEN_13971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13973 = 7'h6b == _myNewVec_20_T_3[6:0] ? myVec_107 : _GEN_13972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13974 = 7'h6c == _myNewVec_20_T_3[6:0] ? myVec_108 : _GEN_13973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13975 = 7'h6d == _myNewVec_20_T_3[6:0] ? myVec_109 : _GEN_13974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13976 = 7'h6e == _myNewVec_20_T_3[6:0] ? myVec_110 : _GEN_13975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13977 = 7'h6f == _myNewVec_20_T_3[6:0] ? myVec_111 : _GEN_13976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13978 = 7'h70 == _myNewVec_20_T_3[6:0] ? myVec_112 : _GEN_13977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13979 = 7'h71 == _myNewVec_20_T_3[6:0] ? myVec_113 : _GEN_13978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13980 = 7'h72 == _myNewVec_20_T_3[6:0] ? myVec_114 : _GEN_13979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13981 = 7'h73 == _myNewVec_20_T_3[6:0] ? myVec_115 : _GEN_13980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13982 = 7'h74 == _myNewVec_20_T_3[6:0] ? myVec_116 : _GEN_13981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13983 = 7'h75 == _myNewVec_20_T_3[6:0] ? myVec_117 : _GEN_13982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13984 = 7'h76 == _myNewVec_20_T_3[6:0] ? myVec_118 : _GEN_13983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13985 = 7'h77 == _myNewVec_20_T_3[6:0] ? myVec_119 : _GEN_13984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13986 = 7'h78 == _myNewVec_20_T_3[6:0] ? myVec_120 : _GEN_13985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13987 = 7'h79 == _myNewVec_20_T_3[6:0] ? myVec_121 : _GEN_13986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13988 = 7'h7a == _myNewVec_20_T_3[6:0] ? myVec_122 : _GEN_13987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13989 = 7'h7b == _myNewVec_20_T_3[6:0] ? myVec_123 : _GEN_13988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13990 = 7'h7c == _myNewVec_20_T_3[6:0] ? myVec_124 : _GEN_13989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13991 = 7'h7d == _myNewVec_20_T_3[6:0] ? myVec_125 : _GEN_13990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13992 = 7'h7e == _myNewVec_20_T_3[6:0] ? myVec_126 : _GEN_13991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_20 = 7'h7f == _myNewVec_20_T_3[6:0] ? myVec_127 : _GEN_13992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_19_T_3 = _myNewVec_127_T_1 + 16'h6c; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_13995 = 7'h1 == _myNewVec_19_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13996 = 7'h2 == _myNewVec_19_T_3[6:0] ? myVec_2 : _GEN_13995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13997 = 7'h3 == _myNewVec_19_T_3[6:0] ? myVec_3 : _GEN_13996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13998 = 7'h4 == _myNewVec_19_T_3[6:0] ? myVec_4 : _GEN_13997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_13999 = 7'h5 == _myNewVec_19_T_3[6:0] ? myVec_5 : _GEN_13998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14000 = 7'h6 == _myNewVec_19_T_3[6:0] ? myVec_6 : _GEN_13999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14001 = 7'h7 == _myNewVec_19_T_3[6:0] ? myVec_7 : _GEN_14000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14002 = 7'h8 == _myNewVec_19_T_3[6:0] ? myVec_8 : _GEN_14001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14003 = 7'h9 == _myNewVec_19_T_3[6:0] ? myVec_9 : _GEN_14002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14004 = 7'ha == _myNewVec_19_T_3[6:0] ? myVec_10 : _GEN_14003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14005 = 7'hb == _myNewVec_19_T_3[6:0] ? myVec_11 : _GEN_14004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14006 = 7'hc == _myNewVec_19_T_3[6:0] ? myVec_12 : _GEN_14005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14007 = 7'hd == _myNewVec_19_T_3[6:0] ? myVec_13 : _GEN_14006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14008 = 7'he == _myNewVec_19_T_3[6:0] ? myVec_14 : _GEN_14007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14009 = 7'hf == _myNewVec_19_T_3[6:0] ? myVec_15 : _GEN_14008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14010 = 7'h10 == _myNewVec_19_T_3[6:0] ? myVec_16 : _GEN_14009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14011 = 7'h11 == _myNewVec_19_T_3[6:0] ? myVec_17 : _GEN_14010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14012 = 7'h12 == _myNewVec_19_T_3[6:0] ? myVec_18 : _GEN_14011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14013 = 7'h13 == _myNewVec_19_T_3[6:0] ? myVec_19 : _GEN_14012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14014 = 7'h14 == _myNewVec_19_T_3[6:0] ? myVec_20 : _GEN_14013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14015 = 7'h15 == _myNewVec_19_T_3[6:0] ? myVec_21 : _GEN_14014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14016 = 7'h16 == _myNewVec_19_T_3[6:0] ? myVec_22 : _GEN_14015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14017 = 7'h17 == _myNewVec_19_T_3[6:0] ? myVec_23 : _GEN_14016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14018 = 7'h18 == _myNewVec_19_T_3[6:0] ? myVec_24 : _GEN_14017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14019 = 7'h19 == _myNewVec_19_T_3[6:0] ? myVec_25 : _GEN_14018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14020 = 7'h1a == _myNewVec_19_T_3[6:0] ? myVec_26 : _GEN_14019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14021 = 7'h1b == _myNewVec_19_T_3[6:0] ? myVec_27 : _GEN_14020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14022 = 7'h1c == _myNewVec_19_T_3[6:0] ? myVec_28 : _GEN_14021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14023 = 7'h1d == _myNewVec_19_T_3[6:0] ? myVec_29 : _GEN_14022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14024 = 7'h1e == _myNewVec_19_T_3[6:0] ? myVec_30 : _GEN_14023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14025 = 7'h1f == _myNewVec_19_T_3[6:0] ? myVec_31 : _GEN_14024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14026 = 7'h20 == _myNewVec_19_T_3[6:0] ? myVec_32 : _GEN_14025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14027 = 7'h21 == _myNewVec_19_T_3[6:0] ? myVec_33 : _GEN_14026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14028 = 7'h22 == _myNewVec_19_T_3[6:0] ? myVec_34 : _GEN_14027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14029 = 7'h23 == _myNewVec_19_T_3[6:0] ? myVec_35 : _GEN_14028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14030 = 7'h24 == _myNewVec_19_T_3[6:0] ? myVec_36 : _GEN_14029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14031 = 7'h25 == _myNewVec_19_T_3[6:0] ? myVec_37 : _GEN_14030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14032 = 7'h26 == _myNewVec_19_T_3[6:0] ? myVec_38 : _GEN_14031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14033 = 7'h27 == _myNewVec_19_T_3[6:0] ? myVec_39 : _GEN_14032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14034 = 7'h28 == _myNewVec_19_T_3[6:0] ? myVec_40 : _GEN_14033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14035 = 7'h29 == _myNewVec_19_T_3[6:0] ? myVec_41 : _GEN_14034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14036 = 7'h2a == _myNewVec_19_T_3[6:0] ? myVec_42 : _GEN_14035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14037 = 7'h2b == _myNewVec_19_T_3[6:0] ? myVec_43 : _GEN_14036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14038 = 7'h2c == _myNewVec_19_T_3[6:0] ? myVec_44 : _GEN_14037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14039 = 7'h2d == _myNewVec_19_T_3[6:0] ? myVec_45 : _GEN_14038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14040 = 7'h2e == _myNewVec_19_T_3[6:0] ? myVec_46 : _GEN_14039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14041 = 7'h2f == _myNewVec_19_T_3[6:0] ? myVec_47 : _GEN_14040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14042 = 7'h30 == _myNewVec_19_T_3[6:0] ? myVec_48 : _GEN_14041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14043 = 7'h31 == _myNewVec_19_T_3[6:0] ? myVec_49 : _GEN_14042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14044 = 7'h32 == _myNewVec_19_T_3[6:0] ? myVec_50 : _GEN_14043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14045 = 7'h33 == _myNewVec_19_T_3[6:0] ? myVec_51 : _GEN_14044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14046 = 7'h34 == _myNewVec_19_T_3[6:0] ? myVec_52 : _GEN_14045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14047 = 7'h35 == _myNewVec_19_T_3[6:0] ? myVec_53 : _GEN_14046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14048 = 7'h36 == _myNewVec_19_T_3[6:0] ? myVec_54 : _GEN_14047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14049 = 7'h37 == _myNewVec_19_T_3[6:0] ? myVec_55 : _GEN_14048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14050 = 7'h38 == _myNewVec_19_T_3[6:0] ? myVec_56 : _GEN_14049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14051 = 7'h39 == _myNewVec_19_T_3[6:0] ? myVec_57 : _GEN_14050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14052 = 7'h3a == _myNewVec_19_T_3[6:0] ? myVec_58 : _GEN_14051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14053 = 7'h3b == _myNewVec_19_T_3[6:0] ? myVec_59 : _GEN_14052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14054 = 7'h3c == _myNewVec_19_T_3[6:0] ? myVec_60 : _GEN_14053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14055 = 7'h3d == _myNewVec_19_T_3[6:0] ? myVec_61 : _GEN_14054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14056 = 7'h3e == _myNewVec_19_T_3[6:0] ? myVec_62 : _GEN_14055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14057 = 7'h3f == _myNewVec_19_T_3[6:0] ? myVec_63 : _GEN_14056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14058 = 7'h40 == _myNewVec_19_T_3[6:0] ? myVec_64 : _GEN_14057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14059 = 7'h41 == _myNewVec_19_T_3[6:0] ? myVec_65 : _GEN_14058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14060 = 7'h42 == _myNewVec_19_T_3[6:0] ? myVec_66 : _GEN_14059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14061 = 7'h43 == _myNewVec_19_T_3[6:0] ? myVec_67 : _GEN_14060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14062 = 7'h44 == _myNewVec_19_T_3[6:0] ? myVec_68 : _GEN_14061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14063 = 7'h45 == _myNewVec_19_T_3[6:0] ? myVec_69 : _GEN_14062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14064 = 7'h46 == _myNewVec_19_T_3[6:0] ? myVec_70 : _GEN_14063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14065 = 7'h47 == _myNewVec_19_T_3[6:0] ? myVec_71 : _GEN_14064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14066 = 7'h48 == _myNewVec_19_T_3[6:0] ? myVec_72 : _GEN_14065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14067 = 7'h49 == _myNewVec_19_T_3[6:0] ? myVec_73 : _GEN_14066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14068 = 7'h4a == _myNewVec_19_T_3[6:0] ? myVec_74 : _GEN_14067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14069 = 7'h4b == _myNewVec_19_T_3[6:0] ? myVec_75 : _GEN_14068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14070 = 7'h4c == _myNewVec_19_T_3[6:0] ? myVec_76 : _GEN_14069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14071 = 7'h4d == _myNewVec_19_T_3[6:0] ? myVec_77 : _GEN_14070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14072 = 7'h4e == _myNewVec_19_T_3[6:0] ? myVec_78 : _GEN_14071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14073 = 7'h4f == _myNewVec_19_T_3[6:0] ? myVec_79 : _GEN_14072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14074 = 7'h50 == _myNewVec_19_T_3[6:0] ? myVec_80 : _GEN_14073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14075 = 7'h51 == _myNewVec_19_T_3[6:0] ? myVec_81 : _GEN_14074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14076 = 7'h52 == _myNewVec_19_T_3[6:0] ? myVec_82 : _GEN_14075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14077 = 7'h53 == _myNewVec_19_T_3[6:0] ? myVec_83 : _GEN_14076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14078 = 7'h54 == _myNewVec_19_T_3[6:0] ? myVec_84 : _GEN_14077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14079 = 7'h55 == _myNewVec_19_T_3[6:0] ? myVec_85 : _GEN_14078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14080 = 7'h56 == _myNewVec_19_T_3[6:0] ? myVec_86 : _GEN_14079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14081 = 7'h57 == _myNewVec_19_T_3[6:0] ? myVec_87 : _GEN_14080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14082 = 7'h58 == _myNewVec_19_T_3[6:0] ? myVec_88 : _GEN_14081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14083 = 7'h59 == _myNewVec_19_T_3[6:0] ? myVec_89 : _GEN_14082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14084 = 7'h5a == _myNewVec_19_T_3[6:0] ? myVec_90 : _GEN_14083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14085 = 7'h5b == _myNewVec_19_T_3[6:0] ? myVec_91 : _GEN_14084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14086 = 7'h5c == _myNewVec_19_T_3[6:0] ? myVec_92 : _GEN_14085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14087 = 7'h5d == _myNewVec_19_T_3[6:0] ? myVec_93 : _GEN_14086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14088 = 7'h5e == _myNewVec_19_T_3[6:0] ? myVec_94 : _GEN_14087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14089 = 7'h5f == _myNewVec_19_T_3[6:0] ? myVec_95 : _GEN_14088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14090 = 7'h60 == _myNewVec_19_T_3[6:0] ? myVec_96 : _GEN_14089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14091 = 7'h61 == _myNewVec_19_T_3[6:0] ? myVec_97 : _GEN_14090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14092 = 7'h62 == _myNewVec_19_T_3[6:0] ? myVec_98 : _GEN_14091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14093 = 7'h63 == _myNewVec_19_T_3[6:0] ? myVec_99 : _GEN_14092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14094 = 7'h64 == _myNewVec_19_T_3[6:0] ? myVec_100 : _GEN_14093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14095 = 7'h65 == _myNewVec_19_T_3[6:0] ? myVec_101 : _GEN_14094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14096 = 7'h66 == _myNewVec_19_T_3[6:0] ? myVec_102 : _GEN_14095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14097 = 7'h67 == _myNewVec_19_T_3[6:0] ? myVec_103 : _GEN_14096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14098 = 7'h68 == _myNewVec_19_T_3[6:0] ? myVec_104 : _GEN_14097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14099 = 7'h69 == _myNewVec_19_T_3[6:0] ? myVec_105 : _GEN_14098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14100 = 7'h6a == _myNewVec_19_T_3[6:0] ? myVec_106 : _GEN_14099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14101 = 7'h6b == _myNewVec_19_T_3[6:0] ? myVec_107 : _GEN_14100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14102 = 7'h6c == _myNewVec_19_T_3[6:0] ? myVec_108 : _GEN_14101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14103 = 7'h6d == _myNewVec_19_T_3[6:0] ? myVec_109 : _GEN_14102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14104 = 7'h6e == _myNewVec_19_T_3[6:0] ? myVec_110 : _GEN_14103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14105 = 7'h6f == _myNewVec_19_T_3[6:0] ? myVec_111 : _GEN_14104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14106 = 7'h70 == _myNewVec_19_T_3[6:0] ? myVec_112 : _GEN_14105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14107 = 7'h71 == _myNewVec_19_T_3[6:0] ? myVec_113 : _GEN_14106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14108 = 7'h72 == _myNewVec_19_T_3[6:0] ? myVec_114 : _GEN_14107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14109 = 7'h73 == _myNewVec_19_T_3[6:0] ? myVec_115 : _GEN_14108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14110 = 7'h74 == _myNewVec_19_T_3[6:0] ? myVec_116 : _GEN_14109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14111 = 7'h75 == _myNewVec_19_T_3[6:0] ? myVec_117 : _GEN_14110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14112 = 7'h76 == _myNewVec_19_T_3[6:0] ? myVec_118 : _GEN_14111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14113 = 7'h77 == _myNewVec_19_T_3[6:0] ? myVec_119 : _GEN_14112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14114 = 7'h78 == _myNewVec_19_T_3[6:0] ? myVec_120 : _GEN_14113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14115 = 7'h79 == _myNewVec_19_T_3[6:0] ? myVec_121 : _GEN_14114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14116 = 7'h7a == _myNewVec_19_T_3[6:0] ? myVec_122 : _GEN_14115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14117 = 7'h7b == _myNewVec_19_T_3[6:0] ? myVec_123 : _GEN_14116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14118 = 7'h7c == _myNewVec_19_T_3[6:0] ? myVec_124 : _GEN_14117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14119 = 7'h7d == _myNewVec_19_T_3[6:0] ? myVec_125 : _GEN_14118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14120 = 7'h7e == _myNewVec_19_T_3[6:0] ? myVec_126 : _GEN_14119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_19 = 7'h7f == _myNewVec_19_T_3[6:0] ? myVec_127 : _GEN_14120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_18_T_3 = _myNewVec_127_T_1 + 16'h6d; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_14123 = 7'h1 == _myNewVec_18_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14124 = 7'h2 == _myNewVec_18_T_3[6:0] ? myVec_2 : _GEN_14123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14125 = 7'h3 == _myNewVec_18_T_3[6:0] ? myVec_3 : _GEN_14124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14126 = 7'h4 == _myNewVec_18_T_3[6:0] ? myVec_4 : _GEN_14125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14127 = 7'h5 == _myNewVec_18_T_3[6:0] ? myVec_5 : _GEN_14126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14128 = 7'h6 == _myNewVec_18_T_3[6:0] ? myVec_6 : _GEN_14127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14129 = 7'h7 == _myNewVec_18_T_3[6:0] ? myVec_7 : _GEN_14128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14130 = 7'h8 == _myNewVec_18_T_3[6:0] ? myVec_8 : _GEN_14129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14131 = 7'h9 == _myNewVec_18_T_3[6:0] ? myVec_9 : _GEN_14130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14132 = 7'ha == _myNewVec_18_T_3[6:0] ? myVec_10 : _GEN_14131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14133 = 7'hb == _myNewVec_18_T_3[6:0] ? myVec_11 : _GEN_14132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14134 = 7'hc == _myNewVec_18_T_3[6:0] ? myVec_12 : _GEN_14133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14135 = 7'hd == _myNewVec_18_T_3[6:0] ? myVec_13 : _GEN_14134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14136 = 7'he == _myNewVec_18_T_3[6:0] ? myVec_14 : _GEN_14135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14137 = 7'hf == _myNewVec_18_T_3[6:0] ? myVec_15 : _GEN_14136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14138 = 7'h10 == _myNewVec_18_T_3[6:0] ? myVec_16 : _GEN_14137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14139 = 7'h11 == _myNewVec_18_T_3[6:0] ? myVec_17 : _GEN_14138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14140 = 7'h12 == _myNewVec_18_T_3[6:0] ? myVec_18 : _GEN_14139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14141 = 7'h13 == _myNewVec_18_T_3[6:0] ? myVec_19 : _GEN_14140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14142 = 7'h14 == _myNewVec_18_T_3[6:0] ? myVec_20 : _GEN_14141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14143 = 7'h15 == _myNewVec_18_T_3[6:0] ? myVec_21 : _GEN_14142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14144 = 7'h16 == _myNewVec_18_T_3[6:0] ? myVec_22 : _GEN_14143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14145 = 7'h17 == _myNewVec_18_T_3[6:0] ? myVec_23 : _GEN_14144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14146 = 7'h18 == _myNewVec_18_T_3[6:0] ? myVec_24 : _GEN_14145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14147 = 7'h19 == _myNewVec_18_T_3[6:0] ? myVec_25 : _GEN_14146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14148 = 7'h1a == _myNewVec_18_T_3[6:0] ? myVec_26 : _GEN_14147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14149 = 7'h1b == _myNewVec_18_T_3[6:0] ? myVec_27 : _GEN_14148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14150 = 7'h1c == _myNewVec_18_T_3[6:0] ? myVec_28 : _GEN_14149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14151 = 7'h1d == _myNewVec_18_T_3[6:0] ? myVec_29 : _GEN_14150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14152 = 7'h1e == _myNewVec_18_T_3[6:0] ? myVec_30 : _GEN_14151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14153 = 7'h1f == _myNewVec_18_T_3[6:0] ? myVec_31 : _GEN_14152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14154 = 7'h20 == _myNewVec_18_T_3[6:0] ? myVec_32 : _GEN_14153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14155 = 7'h21 == _myNewVec_18_T_3[6:0] ? myVec_33 : _GEN_14154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14156 = 7'h22 == _myNewVec_18_T_3[6:0] ? myVec_34 : _GEN_14155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14157 = 7'h23 == _myNewVec_18_T_3[6:0] ? myVec_35 : _GEN_14156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14158 = 7'h24 == _myNewVec_18_T_3[6:0] ? myVec_36 : _GEN_14157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14159 = 7'h25 == _myNewVec_18_T_3[6:0] ? myVec_37 : _GEN_14158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14160 = 7'h26 == _myNewVec_18_T_3[6:0] ? myVec_38 : _GEN_14159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14161 = 7'h27 == _myNewVec_18_T_3[6:0] ? myVec_39 : _GEN_14160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14162 = 7'h28 == _myNewVec_18_T_3[6:0] ? myVec_40 : _GEN_14161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14163 = 7'h29 == _myNewVec_18_T_3[6:0] ? myVec_41 : _GEN_14162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14164 = 7'h2a == _myNewVec_18_T_3[6:0] ? myVec_42 : _GEN_14163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14165 = 7'h2b == _myNewVec_18_T_3[6:0] ? myVec_43 : _GEN_14164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14166 = 7'h2c == _myNewVec_18_T_3[6:0] ? myVec_44 : _GEN_14165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14167 = 7'h2d == _myNewVec_18_T_3[6:0] ? myVec_45 : _GEN_14166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14168 = 7'h2e == _myNewVec_18_T_3[6:0] ? myVec_46 : _GEN_14167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14169 = 7'h2f == _myNewVec_18_T_3[6:0] ? myVec_47 : _GEN_14168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14170 = 7'h30 == _myNewVec_18_T_3[6:0] ? myVec_48 : _GEN_14169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14171 = 7'h31 == _myNewVec_18_T_3[6:0] ? myVec_49 : _GEN_14170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14172 = 7'h32 == _myNewVec_18_T_3[6:0] ? myVec_50 : _GEN_14171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14173 = 7'h33 == _myNewVec_18_T_3[6:0] ? myVec_51 : _GEN_14172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14174 = 7'h34 == _myNewVec_18_T_3[6:0] ? myVec_52 : _GEN_14173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14175 = 7'h35 == _myNewVec_18_T_3[6:0] ? myVec_53 : _GEN_14174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14176 = 7'h36 == _myNewVec_18_T_3[6:0] ? myVec_54 : _GEN_14175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14177 = 7'h37 == _myNewVec_18_T_3[6:0] ? myVec_55 : _GEN_14176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14178 = 7'h38 == _myNewVec_18_T_3[6:0] ? myVec_56 : _GEN_14177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14179 = 7'h39 == _myNewVec_18_T_3[6:0] ? myVec_57 : _GEN_14178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14180 = 7'h3a == _myNewVec_18_T_3[6:0] ? myVec_58 : _GEN_14179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14181 = 7'h3b == _myNewVec_18_T_3[6:0] ? myVec_59 : _GEN_14180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14182 = 7'h3c == _myNewVec_18_T_3[6:0] ? myVec_60 : _GEN_14181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14183 = 7'h3d == _myNewVec_18_T_3[6:0] ? myVec_61 : _GEN_14182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14184 = 7'h3e == _myNewVec_18_T_3[6:0] ? myVec_62 : _GEN_14183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14185 = 7'h3f == _myNewVec_18_T_3[6:0] ? myVec_63 : _GEN_14184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14186 = 7'h40 == _myNewVec_18_T_3[6:0] ? myVec_64 : _GEN_14185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14187 = 7'h41 == _myNewVec_18_T_3[6:0] ? myVec_65 : _GEN_14186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14188 = 7'h42 == _myNewVec_18_T_3[6:0] ? myVec_66 : _GEN_14187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14189 = 7'h43 == _myNewVec_18_T_3[6:0] ? myVec_67 : _GEN_14188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14190 = 7'h44 == _myNewVec_18_T_3[6:0] ? myVec_68 : _GEN_14189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14191 = 7'h45 == _myNewVec_18_T_3[6:0] ? myVec_69 : _GEN_14190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14192 = 7'h46 == _myNewVec_18_T_3[6:0] ? myVec_70 : _GEN_14191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14193 = 7'h47 == _myNewVec_18_T_3[6:0] ? myVec_71 : _GEN_14192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14194 = 7'h48 == _myNewVec_18_T_3[6:0] ? myVec_72 : _GEN_14193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14195 = 7'h49 == _myNewVec_18_T_3[6:0] ? myVec_73 : _GEN_14194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14196 = 7'h4a == _myNewVec_18_T_3[6:0] ? myVec_74 : _GEN_14195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14197 = 7'h4b == _myNewVec_18_T_3[6:0] ? myVec_75 : _GEN_14196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14198 = 7'h4c == _myNewVec_18_T_3[6:0] ? myVec_76 : _GEN_14197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14199 = 7'h4d == _myNewVec_18_T_3[6:0] ? myVec_77 : _GEN_14198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14200 = 7'h4e == _myNewVec_18_T_3[6:0] ? myVec_78 : _GEN_14199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14201 = 7'h4f == _myNewVec_18_T_3[6:0] ? myVec_79 : _GEN_14200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14202 = 7'h50 == _myNewVec_18_T_3[6:0] ? myVec_80 : _GEN_14201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14203 = 7'h51 == _myNewVec_18_T_3[6:0] ? myVec_81 : _GEN_14202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14204 = 7'h52 == _myNewVec_18_T_3[6:0] ? myVec_82 : _GEN_14203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14205 = 7'h53 == _myNewVec_18_T_3[6:0] ? myVec_83 : _GEN_14204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14206 = 7'h54 == _myNewVec_18_T_3[6:0] ? myVec_84 : _GEN_14205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14207 = 7'h55 == _myNewVec_18_T_3[6:0] ? myVec_85 : _GEN_14206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14208 = 7'h56 == _myNewVec_18_T_3[6:0] ? myVec_86 : _GEN_14207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14209 = 7'h57 == _myNewVec_18_T_3[6:0] ? myVec_87 : _GEN_14208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14210 = 7'h58 == _myNewVec_18_T_3[6:0] ? myVec_88 : _GEN_14209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14211 = 7'h59 == _myNewVec_18_T_3[6:0] ? myVec_89 : _GEN_14210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14212 = 7'h5a == _myNewVec_18_T_3[6:0] ? myVec_90 : _GEN_14211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14213 = 7'h5b == _myNewVec_18_T_3[6:0] ? myVec_91 : _GEN_14212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14214 = 7'h5c == _myNewVec_18_T_3[6:0] ? myVec_92 : _GEN_14213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14215 = 7'h5d == _myNewVec_18_T_3[6:0] ? myVec_93 : _GEN_14214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14216 = 7'h5e == _myNewVec_18_T_3[6:0] ? myVec_94 : _GEN_14215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14217 = 7'h5f == _myNewVec_18_T_3[6:0] ? myVec_95 : _GEN_14216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14218 = 7'h60 == _myNewVec_18_T_3[6:0] ? myVec_96 : _GEN_14217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14219 = 7'h61 == _myNewVec_18_T_3[6:0] ? myVec_97 : _GEN_14218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14220 = 7'h62 == _myNewVec_18_T_3[6:0] ? myVec_98 : _GEN_14219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14221 = 7'h63 == _myNewVec_18_T_3[6:0] ? myVec_99 : _GEN_14220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14222 = 7'h64 == _myNewVec_18_T_3[6:0] ? myVec_100 : _GEN_14221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14223 = 7'h65 == _myNewVec_18_T_3[6:0] ? myVec_101 : _GEN_14222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14224 = 7'h66 == _myNewVec_18_T_3[6:0] ? myVec_102 : _GEN_14223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14225 = 7'h67 == _myNewVec_18_T_3[6:0] ? myVec_103 : _GEN_14224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14226 = 7'h68 == _myNewVec_18_T_3[6:0] ? myVec_104 : _GEN_14225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14227 = 7'h69 == _myNewVec_18_T_3[6:0] ? myVec_105 : _GEN_14226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14228 = 7'h6a == _myNewVec_18_T_3[6:0] ? myVec_106 : _GEN_14227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14229 = 7'h6b == _myNewVec_18_T_3[6:0] ? myVec_107 : _GEN_14228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14230 = 7'h6c == _myNewVec_18_T_3[6:0] ? myVec_108 : _GEN_14229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14231 = 7'h6d == _myNewVec_18_T_3[6:0] ? myVec_109 : _GEN_14230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14232 = 7'h6e == _myNewVec_18_T_3[6:0] ? myVec_110 : _GEN_14231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14233 = 7'h6f == _myNewVec_18_T_3[6:0] ? myVec_111 : _GEN_14232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14234 = 7'h70 == _myNewVec_18_T_3[6:0] ? myVec_112 : _GEN_14233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14235 = 7'h71 == _myNewVec_18_T_3[6:0] ? myVec_113 : _GEN_14234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14236 = 7'h72 == _myNewVec_18_T_3[6:0] ? myVec_114 : _GEN_14235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14237 = 7'h73 == _myNewVec_18_T_3[6:0] ? myVec_115 : _GEN_14236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14238 = 7'h74 == _myNewVec_18_T_3[6:0] ? myVec_116 : _GEN_14237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14239 = 7'h75 == _myNewVec_18_T_3[6:0] ? myVec_117 : _GEN_14238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14240 = 7'h76 == _myNewVec_18_T_3[6:0] ? myVec_118 : _GEN_14239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14241 = 7'h77 == _myNewVec_18_T_3[6:0] ? myVec_119 : _GEN_14240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14242 = 7'h78 == _myNewVec_18_T_3[6:0] ? myVec_120 : _GEN_14241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14243 = 7'h79 == _myNewVec_18_T_3[6:0] ? myVec_121 : _GEN_14242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14244 = 7'h7a == _myNewVec_18_T_3[6:0] ? myVec_122 : _GEN_14243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14245 = 7'h7b == _myNewVec_18_T_3[6:0] ? myVec_123 : _GEN_14244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14246 = 7'h7c == _myNewVec_18_T_3[6:0] ? myVec_124 : _GEN_14245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14247 = 7'h7d == _myNewVec_18_T_3[6:0] ? myVec_125 : _GEN_14246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14248 = 7'h7e == _myNewVec_18_T_3[6:0] ? myVec_126 : _GEN_14247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_18 = 7'h7f == _myNewVec_18_T_3[6:0] ? myVec_127 : _GEN_14248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_17_T_3 = _myNewVec_127_T_1 + 16'h6e; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_14251 = 7'h1 == _myNewVec_17_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14252 = 7'h2 == _myNewVec_17_T_3[6:0] ? myVec_2 : _GEN_14251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14253 = 7'h3 == _myNewVec_17_T_3[6:0] ? myVec_3 : _GEN_14252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14254 = 7'h4 == _myNewVec_17_T_3[6:0] ? myVec_4 : _GEN_14253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14255 = 7'h5 == _myNewVec_17_T_3[6:0] ? myVec_5 : _GEN_14254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14256 = 7'h6 == _myNewVec_17_T_3[6:0] ? myVec_6 : _GEN_14255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14257 = 7'h7 == _myNewVec_17_T_3[6:0] ? myVec_7 : _GEN_14256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14258 = 7'h8 == _myNewVec_17_T_3[6:0] ? myVec_8 : _GEN_14257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14259 = 7'h9 == _myNewVec_17_T_3[6:0] ? myVec_9 : _GEN_14258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14260 = 7'ha == _myNewVec_17_T_3[6:0] ? myVec_10 : _GEN_14259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14261 = 7'hb == _myNewVec_17_T_3[6:0] ? myVec_11 : _GEN_14260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14262 = 7'hc == _myNewVec_17_T_3[6:0] ? myVec_12 : _GEN_14261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14263 = 7'hd == _myNewVec_17_T_3[6:0] ? myVec_13 : _GEN_14262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14264 = 7'he == _myNewVec_17_T_3[6:0] ? myVec_14 : _GEN_14263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14265 = 7'hf == _myNewVec_17_T_3[6:0] ? myVec_15 : _GEN_14264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14266 = 7'h10 == _myNewVec_17_T_3[6:0] ? myVec_16 : _GEN_14265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14267 = 7'h11 == _myNewVec_17_T_3[6:0] ? myVec_17 : _GEN_14266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14268 = 7'h12 == _myNewVec_17_T_3[6:0] ? myVec_18 : _GEN_14267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14269 = 7'h13 == _myNewVec_17_T_3[6:0] ? myVec_19 : _GEN_14268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14270 = 7'h14 == _myNewVec_17_T_3[6:0] ? myVec_20 : _GEN_14269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14271 = 7'h15 == _myNewVec_17_T_3[6:0] ? myVec_21 : _GEN_14270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14272 = 7'h16 == _myNewVec_17_T_3[6:0] ? myVec_22 : _GEN_14271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14273 = 7'h17 == _myNewVec_17_T_3[6:0] ? myVec_23 : _GEN_14272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14274 = 7'h18 == _myNewVec_17_T_3[6:0] ? myVec_24 : _GEN_14273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14275 = 7'h19 == _myNewVec_17_T_3[6:0] ? myVec_25 : _GEN_14274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14276 = 7'h1a == _myNewVec_17_T_3[6:0] ? myVec_26 : _GEN_14275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14277 = 7'h1b == _myNewVec_17_T_3[6:0] ? myVec_27 : _GEN_14276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14278 = 7'h1c == _myNewVec_17_T_3[6:0] ? myVec_28 : _GEN_14277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14279 = 7'h1d == _myNewVec_17_T_3[6:0] ? myVec_29 : _GEN_14278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14280 = 7'h1e == _myNewVec_17_T_3[6:0] ? myVec_30 : _GEN_14279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14281 = 7'h1f == _myNewVec_17_T_3[6:0] ? myVec_31 : _GEN_14280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14282 = 7'h20 == _myNewVec_17_T_3[6:0] ? myVec_32 : _GEN_14281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14283 = 7'h21 == _myNewVec_17_T_3[6:0] ? myVec_33 : _GEN_14282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14284 = 7'h22 == _myNewVec_17_T_3[6:0] ? myVec_34 : _GEN_14283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14285 = 7'h23 == _myNewVec_17_T_3[6:0] ? myVec_35 : _GEN_14284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14286 = 7'h24 == _myNewVec_17_T_3[6:0] ? myVec_36 : _GEN_14285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14287 = 7'h25 == _myNewVec_17_T_3[6:0] ? myVec_37 : _GEN_14286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14288 = 7'h26 == _myNewVec_17_T_3[6:0] ? myVec_38 : _GEN_14287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14289 = 7'h27 == _myNewVec_17_T_3[6:0] ? myVec_39 : _GEN_14288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14290 = 7'h28 == _myNewVec_17_T_3[6:0] ? myVec_40 : _GEN_14289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14291 = 7'h29 == _myNewVec_17_T_3[6:0] ? myVec_41 : _GEN_14290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14292 = 7'h2a == _myNewVec_17_T_3[6:0] ? myVec_42 : _GEN_14291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14293 = 7'h2b == _myNewVec_17_T_3[6:0] ? myVec_43 : _GEN_14292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14294 = 7'h2c == _myNewVec_17_T_3[6:0] ? myVec_44 : _GEN_14293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14295 = 7'h2d == _myNewVec_17_T_3[6:0] ? myVec_45 : _GEN_14294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14296 = 7'h2e == _myNewVec_17_T_3[6:0] ? myVec_46 : _GEN_14295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14297 = 7'h2f == _myNewVec_17_T_3[6:0] ? myVec_47 : _GEN_14296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14298 = 7'h30 == _myNewVec_17_T_3[6:0] ? myVec_48 : _GEN_14297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14299 = 7'h31 == _myNewVec_17_T_3[6:0] ? myVec_49 : _GEN_14298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14300 = 7'h32 == _myNewVec_17_T_3[6:0] ? myVec_50 : _GEN_14299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14301 = 7'h33 == _myNewVec_17_T_3[6:0] ? myVec_51 : _GEN_14300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14302 = 7'h34 == _myNewVec_17_T_3[6:0] ? myVec_52 : _GEN_14301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14303 = 7'h35 == _myNewVec_17_T_3[6:0] ? myVec_53 : _GEN_14302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14304 = 7'h36 == _myNewVec_17_T_3[6:0] ? myVec_54 : _GEN_14303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14305 = 7'h37 == _myNewVec_17_T_3[6:0] ? myVec_55 : _GEN_14304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14306 = 7'h38 == _myNewVec_17_T_3[6:0] ? myVec_56 : _GEN_14305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14307 = 7'h39 == _myNewVec_17_T_3[6:0] ? myVec_57 : _GEN_14306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14308 = 7'h3a == _myNewVec_17_T_3[6:0] ? myVec_58 : _GEN_14307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14309 = 7'h3b == _myNewVec_17_T_3[6:0] ? myVec_59 : _GEN_14308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14310 = 7'h3c == _myNewVec_17_T_3[6:0] ? myVec_60 : _GEN_14309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14311 = 7'h3d == _myNewVec_17_T_3[6:0] ? myVec_61 : _GEN_14310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14312 = 7'h3e == _myNewVec_17_T_3[6:0] ? myVec_62 : _GEN_14311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14313 = 7'h3f == _myNewVec_17_T_3[6:0] ? myVec_63 : _GEN_14312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14314 = 7'h40 == _myNewVec_17_T_3[6:0] ? myVec_64 : _GEN_14313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14315 = 7'h41 == _myNewVec_17_T_3[6:0] ? myVec_65 : _GEN_14314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14316 = 7'h42 == _myNewVec_17_T_3[6:0] ? myVec_66 : _GEN_14315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14317 = 7'h43 == _myNewVec_17_T_3[6:0] ? myVec_67 : _GEN_14316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14318 = 7'h44 == _myNewVec_17_T_3[6:0] ? myVec_68 : _GEN_14317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14319 = 7'h45 == _myNewVec_17_T_3[6:0] ? myVec_69 : _GEN_14318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14320 = 7'h46 == _myNewVec_17_T_3[6:0] ? myVec_70 : _GEN_14319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14321 = 7'h47 == _myNewVec_17_T_3[6:0] ? myVec_71 : _GEN_14320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14322 = 7'h48 == _myNewVec_17_T_3[6:0] ? myVec_72 : _GEN_14321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14323 = 7'h49 == _myNewVec_17_T_3[6:0] ? myVec_73 : _GEN_14322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14324 = 7'h4a == _myNewVec_17_T_3[6:0] ? myVec_74 : _GEN_14323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14325 = 7'h4b == _myNewVec_17_T_3[6:0] ? myVec_75 : _GEN_14324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14326 = 7'h4c == _myNewVec_17_T_3[6:0] ? myVec_76 : _GEN_14325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14327 = 7'h4d == _myNewVec_17_T_3[6:0] ? myVec_77 : _GEN_14326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14328 = 7'h4e == _myNewVec_17_T_3[6:0] ? myVec_78 : _GEN_14327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14329 = 7'h4f == _myNewVec_17_T_3[6:0] ? myVec_79 : _GEN_14328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14330 = 7'h50 == _myNewVec_17_T_3[6:0] ? myVec_80 : _GEN_14329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14331 = 7'h51 == _myNewVec_17_T_3[6:0] ? myVec_81 : _GEN_14330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14332 = 7'h52 == _myNewVec_17_T_3[6:0] ? myVec_82 : _GEN_14331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14333 = 7'h53 == _myNewVec_17_T_3[6:0] ? myVec_83 : _GEN_14332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14334 = 7'h54 == _myNewVec_17_T_3[6:0] ? myVec_84 : _GEN_14333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14335 = 7'h55 == _myNewVec_17_T_3[6:0] ? myVec_85 : _GEN_14334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14336 = 7'h56 == _myNewVec_17_T_3[6:0] ? myVec_86 : _GEN_14335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14337 = 7'h57 == _myNewVec_17_T_3[6:0] ? myVec_87 : _GEN_14336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14338 = 7'h58 == _myNewVec_17_T_3[6:0] ? myVec_88 : _GEN_14337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14339 = 7'h59 == _myNewVec_17_T_3[6:0] ? myVec_89 : _GEN_14338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14340 = 7'h5a == _myNewVec_17_T_3[6:0] ? myVec_90 : _GEN_14339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14341 = 7'h5b == _myNewVec_17_T_3[6:0] ? myVec_91 : _GEN_14340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14342 = 7'h5c == _myNewVec_17_T_3[6:0] ? myVec_92 : _GEN_14341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14343 = 7'h5d == _myNewVec_17_T_3[6:0] ? myVec_93 : _GEN_14342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14344 = 7'h5e == _myNewVec_17_T_3[6:0] ? myVec_94 : _GEN_14343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14345 = 7'h5f == _myNewVec_17_T_3[6:0] ? myVec_95 : _GEN_14344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14346 = 7'h60 == _myNewVec_17_T_3[6:0] ? myVec_96 : _GEN_14345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14347 = 7'h61 == _myNewVec_17_T_3[6:0] ? myVec_97 : _GEN_14346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14348 = 7'h62 == _myNewVec_17_T_3[6:0] ? myVec_98 : _GEN_14347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14349 = 7'h63 == _myNewVec_17_T_3[6:0] ? myVec_99 : _GEN_14348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14350 = 7'h64 == _myNewVec_17_T_3[6:0] ? myVec_100 : _GEN_14349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14351 = 7'h65 == _myNewVec_17_T_3[6:0] ? myVec_101 : _GEN_14350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14352 = 7'h66 == _myNewVec_17_T_3[6:0] ? myVec_102 : _GEN_14351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14353 = 7'h67 == _myNewVec_17_T_3[6:0] ? myVec_103 : _GEN_14352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14354 = 7'h68 == _myNewVec_17_T_3[6:0] ? myVec_104 : _GEN_14353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14355 = 7'h69 == _myNewVec_17_T_3[6:0] ? myVec_105 : _GEN_14354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14356 = 7'h6a == _myNewVec_17_T_3[6:0] ? myVec_106 : _GEN_14355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14357 = 7'h6b == _myNewVec_17_T_3[6:0] ? myVec_107 : _GEN_14356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14358 = 7'h6c == _myNewVec_17_T_3[6:0] ? myVec_108 : _GEN_14357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14359 = 7'h6d == _myNewVec_17_T_3[6:0] ? myVec_109 : _GEN_14358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14360 = 7'h6e == _myNewVec_17_T_3[6:0] ? myVec_110 : _GEN_14359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14361 = 7'h6f == _myNewVec_17_T_3[6:0] ? myVec_111 : _GEN_14360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14362 = 7'h70 == _myNewVec_17_T_3[6:0] ? myVec_112 : _GEN_14361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14363 = 7'h71 == _myNewVec_17_T_3[6:0] ? myVec_113 : _GEN_14362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14364 = 7'h72 == _myNewVec_17_T_3[6:0] ? myVec_114 : _GEN_14363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14365 = 7'h73 == _myNewVec_17_T_3[6:0] ? myVec_115 : _GEN_14364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14366 = 7'h74 == _myNewVec_17_T_3[6:0] ? myVec_116 : _GEN_14365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14367 = 7'h75 == _myNewVec_17_T_3[6:0] ? myVec_117 : _GEN_14366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14368 = 7'h76 == _myNewVec_17_T_3[6:0] ? myVec_118 : _GEN_14367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14369 = 7'h77 == _myNewVec_17_T_3[6:0] ? myVec_119 : _GEN_14368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14370 = 7'h78 == _myNewVec_17_T_3[6:0] ? myVec_120 : _GEN_14369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14371 = 7'h79 == _myNewVec_17_T_3[6:0] ? myVec_121 : _GEN_14370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14372 = 7'h7a == _myNewVec_17_T_3[6:0] ? myVec_122 : _GEN_14371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14373 = 7'h7b == _myNewVec_17_T_3[6:0] ? myVec_123 : _GEN_14372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14374 = 7'h7c == _myNewVec_17_T_3[6:0] ? myVec_124 : _GEN_14373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14375 = 7'h7d == _myNewVec_17_T_3[6:0] ? myVec_125 : _GEN_14374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14376 = 7'h7e == _myNewVec_17_T_3[6:0] ? myVec_126 : _GEN_14375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_17 = 7'h7f == _myNewVec_17_T_3[6:0] ? myVec_127 : _GEN_14376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_16_T_3 = _myNewVec_127_T_1 + 16'h6f; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_14379 = 7'h1 == _myNewVec_16_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14380 = 7'h2 == _myNewVec_16_T_3[6:0] ? myVec_2 : _GEN_14379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14381 = 7'h3 == _myNewVec_16_T_3[6:0] ? myVec_3 : _GEN_14380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14382 = 7'h4 == _myNewVec_16_T_3[6:0] ? myVec_4 : _GEN_14381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14383 = 7'h5 == _myNewVec_16_T_3[6:0] ? myVec_5 : _GEN_14382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14384 = 7'h6 == _myNewVec_16_T_3[6:0] ? myVec_6 : _GEN_14383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14385 = 7'h7 == _myNewVec_16_T_3[6:0] ? myVec_7 : _GEN_14384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14386 = 7'h8 == _myNewVec_16_T_3[6:0] ? myVec_8 : _GEN_14385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14387 = 7'h9 == _myNewVec_16_T_3[6:0] ? myVec_9 : _GEN_14386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14388 = 7'ha == _myNewVec_16_T_3[6:0] ? myVec_10 : _GEN_14387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14389 = 7'hb == _myNewVec_16_T_3[6:0] ? myVec_11 : _GEN_14388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14390 = 7'hc == _myNewVec_16_T_3[6:0] ? myVec_12 : _GEN_14389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14391 = 7'hd == _myNewVec_16_T_3[6:0] ? myVec_13 : _GEN_14390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14392 = 7'he == _myNewVec_16_T_3[6:0] ? myVec_14 : _GEN_14391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14393 = 7'hf == _myNewVec_16_T_3[6:0] ? myVec_15 : _GEN_14392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14394 = 7'h10 == _myNewVec_16_T_3[6:0] ? myVec_16 : _GEN_14393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14395 = 7'h11 == _myNewVec_16_T_3[6:0] ? myVec_17 : _GEN_14394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14396 = 7'h12 == _myNewVec_16_T_3[6:0] ? myVec_18 : _GEN_14395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14397 = 7'h13 == _myNewVec_16_T_3[6:0] ? myVec_19 : _GEN_14396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14398 = 7'h14 == _myNewVec_16_T_3[6:0] ? myVec_20 : _GEN_14397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14399 = 7'h15 == _myNewVec_16_T_3[6:0] ? myVec_21 : _GEN_14398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14400 = 7'h16 == _myNewVec_16_T_3[6:0] ? myVec_22 : _GEN_14399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14401 = 7'h17 == _myNewVec_16_T_3[6:0] ? myVec_23 : _GEN_14400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14402 = 7'h18 == _myNewVec_16_T_3[6:0] ? myVec_24 : _GEN_14401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14403 = 7'h19 == _myNewVec_16_T_3[6:0] ? myVec_25 : _GEN_14402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14404 = 7'h1a == _myNewVec_16_T_3[6:0] ? myVec_26 : _GEN_14403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14405 = 7'h1b == _myNewVec_16_T_3[6:0] ? myVec_27 : _GEN_14404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14406 = 7'h1c == _myNewVec_16_T_3[6:0] ? myVec_28 : _GEN_14405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14407 = 7'h1d == _myNewVec_16_T_3[6:0] ? myVec_29 : _GEN_14406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14408 = 7'h1e == _myNewVec_16_T_3[6:0] ? myVec_30 : _GEN_14407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14409 = 7'h1f == _myNewVec_16_T_3[6:0] ? myVec_31 : _GEN_14408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14410 = 7'h20 == _myNewVec_16_T_3[6:0] ? myVec_32 : _GEN_14409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14411 = 7'h21 == _myNewVec_16_T_3[6:0] ? myVec_33 : _GEN_14410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14412 = 7'h22 == _myNewVec_16_T_3[6:0] ? myVec_34 : _GEN_14411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14413 = 7'h23 == _myNewVec_16_T_3[6:0] ? myVec_35 : _GEN_14412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14414 = 7'h24 == _myNewVec_16_T_3[6:0] ? myVec_36 : _GEN_14413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14415 = 7'h25 == _myNewVec_16_T_3[6:0] ? myVec_37 : _GEN_14414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14416 = 7'h26 == _myNewVec_16_T_3[6:0] ? myVec_38 : _GEN_14415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14417 = 7'h27 == _myNewVec_16_T_3[6:0] ? myVec_39 : _GEN_14416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14418 = 7'h28 == _myNewVec_16_T_3[6:0] ? myVec_40 : _GEN_14417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14419 = 7'h29 == _myNewVec_16_T_3[6:0] ? myVec_41 : _GEN_14418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14420 = 7'h2a == _myNewVec_16_T_3[6:0] ? myVec_42 : _GEN_14419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14421 = 7'h2b == _myNewVec_16_T_3[6:0] ? myVec_43 : _GEN_14420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14422 = 7'h2c == _myNewVec_16_T_3[6:0] ? myVec_44 : _GEN_14421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14423 = 7'h2d == _myNewVec_16_T_3[6:0] ? myVec_45 : _GEN_14422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14424 = 7'h2e == _myNewVec_16_T_3[6:0] ? myVec_46 : _GEN_14423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14425 = 7'h2f == _myNewVec_16_T_3[6:0] ? myVec_47 : _GEN_14424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14426 = 7'h30 == _myNewVec_16_T_3[6:0] ? myVec_48 : _GEN_14425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14427 = 7'h31 == _myNewVec_16_T_3[6:0] ? myVec_49 : _GEN_14426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14428 = 7'h32 == _myNewVec_16_T_3[6:0] ? myVec_50 : _GEN_14427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14429 = 7'h33 == _myNewVec_16_T_3[6:0] ? myVec_51 : _GEN_14428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14430 = 7'h34 == _myNewVec_16_T_3[6:0] ? myVec_52 : _GEN_14429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14431 = 7'h35 == _myNewVec_16_T_3[6:0] ? myVec_53 : _GEN_14430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14432 = 7'h36 == _myNewVec_16_T_3[6:0] ? myVec_54 : _GEN_14431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14433 = 7'h37 == _myNewVec_16_T_3[6:0] ? myVec_55 : _GEN_14432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14434 = 7'h38 == _myNewVec_16_T_3[6:0] ? myVec_56 : _GEN_14433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14435 = 7'h39 == _myNewVec_16_T_3[6:0] ? myVec_57 : _GEN_14434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14436 = 7'h3a == _myNewVec_16_T_3[6:0] ? myVec_58 : _GEN_14435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14437 = 7'h3b == _myNewVec_16_T_3[6:0] ? myVec_59 : _GEN_14436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14438 = 7'h3c == _myNewVec_16_T_3[6:0] ? myVec_60 : _GEN_14437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14439 = 7'h3d == _myNewVec_16_T_3[6:0] ? myVec_61 : _GEN_14438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14440 = 7'h3e == _myNewVec_16_T_3[6:0] ? myVec_62 : _GEN_14439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14441 = 7'h3f == _myNewVec_16_T_3[6:0] ? myVec_63 : _GEN_14440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14442 = 7'h40 == _myNewVec_16_T_3[6:0] ? myVec_64 : _GEN_14441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14443 = 7'h41 == _myNewVec_16_T_3[6:0] ? myVec_65 : _GEN_14442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14444 = 7'h42 == _myNewVec_16_T_3[6:0] ? myVec_66 : _GEN_14443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14445 = 7'h43 == _myNewVec_16_T_3[6:0] ? myVec_67 : _GEN_14444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14446 = 7'h44 == _myNewVec_16_T_3[6:0] ? myVec_68 : _GEN_14445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14447 = 7'h45 == _myNewVec_16_T_3[6:0] ? myVec_69 : _GEN_14446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14448 = 7'h46 == _myNewVec_16_T_3[6:0] ? myVec_70 : _GEN_14447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14449 = 7'h47 == _myNewVec_16_T_3[6:0] ? myVec_71 : _GEN_14448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14450 = 7'h48 == _myNewVec_16_T_3[6:0] ? myVec_72 : _GEN_14449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14451 = 7'h49 == _myNewVec_16_T_3[6:0] ? myVec_73 : _GEN_14450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14452 = 7'h4a == _myNewVec_16_T_3[6:0] ? myVec_74 : _GEN_14451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14453 = 7'h4b == _myNewVec_16_T_3[6:0] ? myVec_75 : _GEN_14452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14454 = 7'h4c == _myNewVec_16_T_3[6:0] ? myVec_76 : _GEN_14453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14455 = 7'h4d == _myNewVec_16_T_3[6:0] ? myVec_77 : _GEN_14454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14456 = 7'h4e == _myNewVec_16_T_3[6:0] ? myVec_78 : _GEN_14455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14457 = 7'h4f == _myNewVec_16_T_3[6:0] ? myVec_79 : _GEN_14456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14458 = 7'h50 == _myNewVec_16_T_3[6:0] ? myVec_80 : _GEN_14457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14459 = 7'h51 == _myNewVec_16_T_3[6:0] ? myVec_81 : _GEN_14458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14460 = 7'h52 == _myNewVec_16_T_3[6:0] ? myVec_82 : _GEN_14459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14461 = 7'h53 == _myNewVec_16_T_3[6:0] ? myVec_83 : _GEN_14460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14462 = 7'h54 == _myNewVec_16_T_3[6:0] ? myVec_84 : _GEN_14461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14463 = 7'h55 == _myNewVec_16_T_3[6:0] ? myVec_85 : _GEN_14462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14464 = 7'h56 == _myNewVec_16_T_3[6:0] ? myVec_86 : _GEN_14463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14465 = 7'h57 == _myNewVec_16_T_3[6:0] ? myVec_87 : _GEN_14464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14466 = 7'h58 == _myNewVec_16_T_3[6:0] ? myVec_88 : _GEN_14465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14467 = 7'h59 == _myNewVec_16_T_3[6:0] ? myVec_89 : _GEN_14466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14468 = 7'h5a == _myNewVec_16_T_3[6:0] ? myVec_90 : _GEN_14467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14469 = 7'h5b == _myNewVec_16_T_3[6:0] ? myVec_91 : _GEN_14468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14470 = 7'h5c == _myNewVec_16_T_3[6:0] ? myVec_92 : _GEN_14469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14471 = 7'h5d == _myNewVec_16_T_3[6:0] ? myVec_93 : _GEN_14470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14472 = 7'h5e == _myNewVec_16_T_3[6:0] ? myVec_94 : _GEN_14471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14473 = 7'h5f == _myNewVec_16_T_3[6:0] ? myVec_95 : _GEN_14472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14474 = 7'h60 == _myNewVec_16_T_3[6:0] ? myVec_96 : _GEN_14473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14475 = 7'h61 == _myNewVec_16_T_3[6:0] ? myVec_97 : _GEN_14474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14476 = 7'h62 == _myNewVec_16_T_3[6:0] ? myVec_98 : _GEN_14475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14477 = 7'h63 == _myNewVec_16_T_3[6:0] ? myVec_99 : _GEN_14476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14478 = 7'h64 == _myNewVec_16_T_3[6:0] ? myVec_100 : _GEN_14477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14479 = 7'h65 == _myNewVec_16_T_3[6:0] ? myVec_101 : _GEN_14478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14480 = 7'h66 == _myNewVec_16_T_3[6:0] ? myVec_102 : _GEN_14479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14481 = 7'h67 == _myNewVec_16_T_3[6:0] ? myVec_103 : _GEN_14480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14482 = 7'h68 == _myNewVec_16_T_3[6:0] ? myVec_104 : _GEN_14481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14483 = 7'h69 == _myNewVec_16_T_3[6:0] ? myVec_105 : _GEN_14482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14484 = 7'h6a == _myNewVec_16_T_3[6:0] ? myVec_106 : _GEN_14483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14485 = 7'h6b == _myNewVec_16_T_3[6:0] ? myVec_107 : _GEN_14484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14486 = 7'h6c == _myNewVec_16_T_3[6:0] ? myVec_108 : _GEN_14485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14487 = 7'h6d == _myNewVec_16_T_3[6:0] ? myVec_109 : _GEN_14486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14488 = 7'h6e == _myNewVec_16_T_3[6:0] ? myVec_110 : _GEN_14487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14489 = 7'h6f == _myNewVec_16_T_3[6:0] ? myVec_111 : _GEN_14488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14490 = 7'h70 == _myNewVec_16_T_3[6:0] ? myVec_112 : _GEN_14489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14491 = 7'h71 == _myNewVec_16_T_3[6:0] ? myVec_113 : _GEN_14490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14492 = 7'h72 == _myNewVec_16_T_3[6:0] ? myVec_114 : _GEN_14491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14493 = 7'h73 == _myNewVec_16_T_3[6:0] ? myVec_115 : _GEN_14492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14494 = 7'h74 == _myNewVec_16_T_3[6:0] ? myVec_116 : _GEN_14493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14495 = 7'h75 == _myNewVec_16_T_3[6:0] ? myVec_117 : _GEN_14494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14496 = 7'h76 == _myNewVec_16_T_3[6:0] ? myVec_118 : _GEN_14495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14497 = 7'h77 == _myNewVec_16_T_3[6:0] ? myVec_119 : _GEN_14496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14498 = 7'h78 == _myNewVec_16_T_3[6:0] ? myVec_120 : _GEN_14497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14499 = 7'h79 == _myNewVec_16_T_3[6:0] ? myVec_121 : _GEN_14498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14500 = 7'h7a == _myNewVec_16_T_3[6:0] ? myVec_122 : _GEN_14499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14501 = 7'h7b == _myNewVec_16_T_3[6:0] ? myVec_123 : _GEN_14500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14502 = 7'h7c == _myNewVec_16_T_3[6:0] ? myVec_124 : _GEN_14501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14503 = 7'h7d == _myNewVec_16_T_3[6:0] ? myVec_125 : _GEN_14502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14504 = 7'h7e == _myNewVec_16_T_3[6:0] ? myVec_126 : _GEN_14503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_16 = 7'h7f == _myNewVec_16_T_3[6:0] ? myVec_127 : _GEN_14504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [255:0] myNewWire_lo_lo_hi_lo = {myNewVec_23,myNewVec_22,myNewVec_21,myNewVec_20,myNewVec_19,myNewVec_18,
    myNewVec_17,myNewVec_16}; // @[hh_datapath_chisel.scala 238:27]
  wire [15:0] _myNewVec_15_T_3 = _myNewVec_127_T_1 + 16'h70; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_14507 = 7'h1 == _myNewVec_15_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14508 = 7'h2 == _myNewVec_15_T_3[6:0] ? myVec_2 : _GEN_14507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14509 = 7'h3 == _myNewVec_15_T_3[6:0] ? myVec_3 : _GEN_14508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14510 = 7'h4 == _myNewVec_15_T_3[6:0] ? myVec_4 : _GEN_14509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14511 = 7'h5 == _myNewVec_15_T_3[6:0] ? myVec_5 : _GEN_14510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14512 = 7'h6 == _myNewVec_15_T_3[6:0] ? myVec_6 : _GEN_14511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14513 = 7'h7 == _myNewVec_15_T_3[6:0] ? myVec_7 : _GEN_14512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14514 = 7'h8 == _myNewVec_15_T_3[6:0] ? myVec_8 : _GEN_14513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14515 = 7'h9 == _myNewVec_15_T_3[6:0] ? myVec_9 : _GEN_14514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14516 = 7'ha == _myNewVec_15_T_3[6:0] ? myVec_10 : _GEN_14515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14517 = 7'hb == _myNewVec_15_T_3[6:0] ? myVec_11 : _GEN_14516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14518 = 7'hc == _myNewVec_15_T_3[6:0] ? myVec_12 : _GEN_14517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14519 = 7'hd == _myNewVec_15_T_3[6:0] ? myVec_13 : _GEN_14518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14520 = 7'he == _myNewVec_15_T_3[6:0] ? myVec_14 : _GEN_14519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14521 = 7'hf == _myNewVec_15_T_3[6:0] ? myVec_15 : _GEN_14520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14522 = 7'h10 == _myNewVec_15_T_3[6:0] ? myVec_16 : _GEN_14521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14523 = 7'h11 == _myNewVec_15_T_3[6:0] ? myVec_17 : _GEN_14522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14524 = 7'h12 == _myNewVec_15_T_3[6:0] ? myVec_18 : _GEN_14523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14525 = 7'h13 == _myNewVec_15_T_3[6:0] ? myVec_19 : _GEN_14524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14526 = 7'h14 == _myNewVec_15_T_3[6:0] ? myVec_20 : _GEN_14525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14527 = 7'h15 == _myNewVec_15_T_3[6:0] ? myVec_21 : _GEN_14526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14528 = 7'h16 == _myNewVec_15_T_3[6:0] ? myVec_22 : _GEN_14527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14529 = 7'h17 == _myNewVec_15_T_3[6:0] ? myVec_23 : _GEN_14528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14530 = 7'h18 == _myNewVec_15_T_3[6:0] ? myVec_24 : _GEN_14529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14531 = 7'h19 == _myNewVec_15_T_3[6:0] ? myVec_25 : _GEN_14530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14532 = 7'h1a == _myNewVec_15_T_3[6:0] ? myVec_26 : _GEN_14531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14533 = 7'h1b == _myNewVec_15_T_3[6:0] ? myVec_27 : _GEN_14532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14534 = 7'h1c == _myNewVec_15_T_3[6:0] ? myVec_28 : _GEN_14533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14535 = 7'h1d == _myNewVec_15_T_3[6:0] ? myVec_29 : _GEN_14534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14536 = 7'h1e == _myNewVec_15_T_3[6:0] ? myVec_30 : _GEN_14535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14537 = 7'h1f == _myNewVec_15_T_3[6:0] ? myVec_31 : _GEN_14536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14538 = 7'h20 == _myNewVec_15_T_3[6:0] ? myVec_32 : _GEN_14537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14539 = 7'h21 == _myNewVec_15_T_3[6:0] ? myVec_33 : _GEN_14538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14540 = 7'h22 == _myNewVec_15_T_3[6:0] ? myVec_34 : _GEN_14539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14541 = 7'h23 == _myNewVec_15_T_3[6:0] ? myVec_35 : _GEN_14540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14542 = 7'h24 == _myNewVec_15_T_3[6:0] ? myVec_36 : _GEN_14541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14543 = 7'h25 == _myNewVec_15_T_3[6:0] ? myVec_37 : _GEN_14542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14544 = 7'h26 == _myNewVec_15_T_3[6:0] ? myVec_38 : _GEN_14543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14545 = 7'h27 == _myNewVec_15_T_3[6:0] ? myVec_39 : _GEN_14544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14546 = 7'h28 == _myNewVec_15_T_3[6:0] ? myVec_40 : _GEN_14545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14547 = 7'h29 == _myNewVec_15_T_3[6:0] ? myVec_41 : _GEN_14546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14548 = 7'h2a == _myNewVec_15_T_3[6:0] ? myVec_42 : _GEN_14547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14549 = 7'h2b == _myNewVec_15_T_3[6:0] ? myVec_43 : _GEN_14548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14550 = 7'h2c == _myNewVec_15_T_3[6:0] ? myVec_44 : _GEN_14549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14551 = 7'h2d == _myNewVec_15_T_3[6:0] ? myVec_45 : _GEN_14550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14552 = 7'h2e == _myNewVec_15_T_3[6:0] ? myVec_46 : _GEN_14551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14553 = 7'h2f == _myNewVec_15_T_3[6:0] ? myVec_47 : _GEN_14552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14554 = 7'h30 == _myNewVec_15_T_3[6:0] ? myVec_48 : _GEN_14553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14555 = 7'h31 == _myNewVec_15_T_3[6:0] ? myVec_49 : _GEN_14554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14556 = 7'h32 == _myNewVec_15_T_3[6:0] ? myVec_50 : _GEN_14555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14557 = 7'h33 == _myNewVec_15_T_3[6:0] ? myVec_51 : _GEN_14556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14558 = 7'h34 == _myNewVec_15_T_3[6:0] ? myVec_52 : _GEN_14557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14559 = 7'h35 == _myNewVec_15_T_3[6:0] ? myVec_53 : _GEN_14558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14560 = 7'h36 == _myNewVec_15_T_3[6:0] ? myVec_54 : _GEN_14559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14561 = 7'h37 == _myNewVec_15_T_3[6:0] ? myVec_55 : _GEN_14560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14562 = 7'h38 == _myNewVec_15_T_3[6:0] ? myVec_56 : _GEN_14561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14563 = 7'h39 == _myNewVec_15_T_3[6:0] ? myVec_57 : _GEN_14562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14564 = 7'h3a == _myNewVec_15_T_3[6:0] ? myVec_58 : _GEN_14563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14565 = 7'h3b == _myNewVec_15_T_3[6:0] ? myVec_59 : _GEN_14564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14566 = 7'h3c == _myNewVec_15_T_3[6:0] ? myVec_60 : _GEN_14565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14567 = 7'h3d == _myNewVec_15_T_3[6:0] ? myVec_61 : _GEN_14566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14568 = 7'h3e == _myNewVec_15_T_3[6:0] ? myVec_62 : _GEN_14567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14569 = 7'h3f == _myNewVec_15_T_3[6:0] ? myVec_63 : _GEN_14568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14570 = 7'h40 == _myNewVec_15_T_3[6:0] ? myVec_64 : _GEN_14569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14571 = 7'h41 == _myNewVec_15_T_3[6:0] ? myVec_65 : _GEN_14570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14572 = 7'h42 == _myNewVec_15_T_3[6:0] ? myVec_66 : _GEN_14571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14573 = 7'h43 == _myNewVec_15_T_3[6:0] ? myVec_67 : _GEN_14572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14574 = 7'h44 == _myNewVec_15_T_3[6:0] ? myVec_68 : _GEN_14573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14575 = 7'h45 == _myNewVec_15_T_3[6:0] ? myVec_69 : _GEN_14574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14576 = 7'h46 == _myNewVec_15_T_3[6:0] ? myVec_70 : _GEN_14575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14577 = 7'h47 == _myNewVec_15_T_3[6:0] ? myVec_71 : _GEN_14576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14578 = 7'h48 == _myNewVec_15_T_3[6:0] ? myVec_72 : _GEN_14577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14579 = 7'h49 == _myNewVec_15_T_3[6:0] ? myVec_73 : _GEN_14578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14580 = 7'h4a == _myNewVec_15_T_3[6:0] ? myVec_74 : _GEN_14579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14581 = 7'h4b == _myNewVec_15_T_3[6:0] ? myVec_75 : _GEN_14580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14582 = 7'h4c == _myNewVec_15_T_3[6:0] ? myVec_76 : _GEN_14581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14583 = 7'h4d == _myNewVec_15_T_3[6:0] ? myVec_77 : _GEN_14582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14584 = 7'h4e == _myNewVec_15_T_3[6:0] ? myVec_78 : _GEN_14583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14585 = 7'h4f == _myNewVec_15_T_3[6:0] ? myVec_79 : _GEN_14584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14586 = 7'h50 == _myNewVec_15_T_3[6:0] ? myVec_80 : _GEN_14585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14587 = 7'h51 == _myNewVec_15_T_3[6:0] ? myVec_81 : _GEN_14586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14588 = 7'h52 == _myNewVec_15_T_3[6:0] ? myVec_82 : _GEN_14587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14589 = 7'h53 == _myNewVec_15_T_3[6:0] ? myVec_83 : _GEN_14588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14590 = 7'h54 == _myNewVec_15_T_3[6:0] ? myVec_84 : _GEN_14589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14591 = 7'h55 == _myNewVec_15_T_3[6:0] ? myVec_85 : _GEN_14590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14592 = 7'h56 == _myNewVec_15_T_3[6:0] ? myVec_86 : _GEN_14591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14593 = 7'h57 == _myNewVec_15_T_3[6:0] ? myVec_87 : _GEN_14592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14594 = 7'h58 == _myNewVec_15_T_3[6:0] ? myVec_88 : _GEN_14593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14595 = 7'h59 == _myNewVec_15_T_3[6:0] ? myVec_89 : _GEN_14594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14596 = 7'h5a == _myNewVec_15_T_3[6:0] ? myVec_90 : _GEN_14595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14597 = 7'h5b == _myNewVec_15_T_3[6:0] ? myVec_91 : _GEN_14596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14598 = 7'h5c == _myNewVec_15_T_3[6:0] ? myVec_92 : _GEN_14597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14599 = 7'h5d == _myNewVec_15_T_3[6:0] ? myVec_93 : _GEN_14598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14600 = 7'h5e == _myNewVec_15_T_3[6:0] ? myVec_94 : _GEN_14599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14601 = 7'h5f == _myNewVec_15_T_3[6:0] ? myVec_95 : _GEN_14600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14602 = 7'h60 == _myNewVec_15_T_3[6:0] ? myVec_96 : _GEN_14601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14603 = 7'h61 == _myNewVec_15_T_3[6:0] ? myVec_97 : _GEN_14602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14604 = 7'h62 == _myNewVec_15_T_3[6:0] ? myVec_98 : _GEN_14603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14605 = 7'h63 == _myNewVec_15_T_3[6:0] ? myVec_99 : _GEN_14604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14606 = 7'h64 == _myNewVec_15_T_3[6:0] ? myVec_100 : _GEN_14605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14607 = 7'h65 == _myNewVec_15_T_3[6:0] ? myVec_101 : _GEN_14606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14608 = 7'h66 == _myNewVec_15_T_3[6:0] ? myVec_102 : _GEN_14607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14609 = 7'h67 == _myNewVec_15_T_3[6:0] ? myVec_103 : _GEN_14608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14610 = 7'h68 == _myNewVec_15_T_3[6:0] ? myVec_104 : _GEN_14609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14611 = 7'h69 == _myNewVec_15_T_3[6:0] ? myVec_105 : _GEN_14610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14612 = 7'h6a == _myNewVec_15_T_3[6:0] ? myVec_106 : _GEN_14611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14613 = 7'h6b == _myNewVec_15_T_3[6:0] ? myVec_107 : _GEN_14612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14614 = 7'h6c == _myNewVec_15_T_3[6:0] ? myVec_108 : _GEN_14613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14615 = 7'h6d == _myNewVec_15_T_3[6:0] ? myVec_109 : _GEN_14614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14616 = 7'h6e == _myNewVec_15_T_3[6:0] ? myVec_110 : _GEN_14615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14617 = 7'h6f == _myNewVec_15_T_3[6:0] ? myVec_111 : _GEN_14616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14618 = 7'h70 == _myNewVec_15_T_3[6:0] ? myVec_112 : _GEN_14617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14619 = 7'h71 == _myNewVec_15_T_3[6:0] ? myVec_113 : _GEN_14618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14620 = 7'h72 == _myNewVec_15_T_3[6:0] ? myVec_114 : _GEN_14619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14621 = 7'h73 == _myNewVec_15_T_3[6:0] ? myVec_115 : _GEN_14620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14622 = 7'h74 == _myNewVec_15_T_3[6:0] ? myVec_116 : _GEN_14621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14623 = 7'h75 == _myNewVec_15_T_3[6:0] ? myVec_117 : _GEN_14622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14624 = 7'h76 == _myNewVec_15_T_3[6:0] ? myVec_118 : _GEN_14623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14625 = 7'h77 == _myNewVec_15_T_3[6:0] ? myVec_119 : _GEN_14624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14626 = 7'h78 == _myNewVec_15_T_3[6:0] ? myVec_120 : _GEN_14625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14627 = 7'h79 == _myNewVec_15_T_3[6:0] ? myVec_121 : _GEN_14626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14628 = 7'h7a == _myNewVec_15_T_3[6:0] ? myVec_122 : _GEN_14627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14629 = 7'h7b == _myNewVec_15_T_3[6:0] ? myVec_123 : _GEN_14628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14630 = 7'h7c == _myNewVec_15_T_3[6:0] ? myVec_124 : _GEN_14629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14631 = 7'h7d == _myNewVec_15_T_3[6:0] ? myVec_125 : _GEN_14630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14632 = 7'h7e == _myNewVec_15_T_3[6:0] ? myVec_126 : _GEN_14631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_15 = 7'h7f == _myNewVec_15_T_3[6:0] ? myVec_127 : _GEN_14632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_14_T_3 = _myNewVec_127_T_1 + 16'h71; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_14635 = 7'h1 == _myNewVec_14_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14636 = 7'h2 == _myNewVec_14_T_3[6:0] ? myVec_2 : _GEN_14635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14637 = 7'h3 == _myNewVec_14_T_3[6:0] ? myVec_3 : _GEN_14636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14638 = 7'h4 == _myNewVec_14_T_3[6:0] ? myVec_4 : _GEN_14637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14639 = 7'h5 == _myNewVec_14_T_3[6:0] ? myVec_5 : _GEN_14638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14640 = 7'h6 == _myNewVec_14_T_3[6:0] ? myVec_6 : _GEN_14639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14641 = 7'h7 == _myNewVec_14_T_3[6:0] ? myVec_7 : _GEN_14640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14642 = 7'h8 == _myNewVec_14_T_3[6:0] ? myVec_8 : _GEN_14641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14643 = 7'h9 == _myNewVec_14_T_3[6:0] ? myVec_9 : _GEN_14642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14644 = 7'ha == _myNewVec_14_T_3[6:0] ? myVec_10 : _GEN_14643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14645 = 7'hb == _myNewVec_14_T_3[6:0] ? myVec_11 : _GEN_14644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14646 = 7'hc == _myNewVec_14_T_3[6:0] ? myVec_12 : _GEN_14645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14647 = 7'hd == _myNewVec_14_T_3[6:0] ? myVec_13 : _GEN_14646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14648 = 7'he == _myNewVec_14_T_3[6:0] ? myVec_14 : _GEN_14647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14649 = 7'hf == _myNewVec_14_T_3[6:0] ? myVec_15 : _GEN_14648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14650 = 7'h10 == _myNewVec_14_T_3[6:0] ? myVec_16 : _GEN_14649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14651 = 7'h11 == _myNewVec_14_T_3[6:0] ? myVec_17 : _GEN_14650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14652 = 7'h12 == _myNewVec_14_T_3[6:0] ? myVec_18 : _GEN_14651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14653 = 7'h13 == _myNewVec_14_T_3[6:0] ? myVec_19 : _GEN_14652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14654 = 7'h14 == _myNewVec_14_T_3[6:0] ? myVec_20 : _GEN_14653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14655 = 7'h15 == _myNewVec_14_T_3[6:0] ? myVec_21 : _GEN_14654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14656 = 7'h16 == _myNewVec_14_T_3[6:0] ? myVec_22 : _GEN_14655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14657 = 7'h17 == _myNewVec_14_T_3[6:0] ? myVec_23 : _GEN_14656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14658 = 7'h18 == _myNewVec_14_T_3[6:0] ? myVec_24 : _GEN_14657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14659 = 7'h19 == _myNewVec_14_T_3[6:0] ? myVec_25 : _GEN_14658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14660 = 7'h1a == _myNewVec_14_T_3[6:0] ? myVec_26 : _GEN_14659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14661 = 7'h1b == _myNewVec_14_T_3[6:0] ? myVec_27 : _GEN_14660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14662 = 7'h1c == _myNewVec_14_T_3[6:0] ? myVec_28 : _GEN_14661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14663 = 7'h1d == _myNewVec_14_T_3[6:0] ? myVec_29 : _GEN_14662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14664 = 7'h1e == _myNewVec_14_T_3[6:0] ? myVec_30 : _GEN_14663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14665 = 7'h1f == _myNewVec_14_T_3[6:0] ? myVec_31 : _GEN_14664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14666 = 7'h20 == _myNewVec_14_T_3[6:0] ? myVec_32 : _GEN_14665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14667 = 7'h21 == _myNewVec_14_T_3[6:0] ? myVec_33 : _GEN_14666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14668 = 7'h22 == _myNewVec_14_T_3[6:0] ? myVec_34 : _GEN_14667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14669 = 7'h23 == _myNewVec_14_T_3[6:0] ? myVec_35 : _GEN_14668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14670 = 7'h24 == _myNewVec_14_T_3[6:0] ? myVec_36 : _GEN_14669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14671 = 7'h25 == _myNewVec_14_T_3[6:0] ? myVec_37 : _GEN_14670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14672 = 7'h26 == _myNewVec_14_T_3[6:0] ? myVec_38 : _GEN_14671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14673 = 7'h27 == _myNewVec_14_T_3[6:0] ? myVec_39 : _GEN_14672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14674 = 7'h28 == _myNewVec_14_T_3[6:0] ? myVec_40 : _GEN_14673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14675 = 7'h29 == _myNewVec_14_T_3[6:0] ? myVec_41 : _GEN_14674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14676 = 7'h2a == _myNewVec_14_T_3[6:0] ? myVec_42 : _GEN_14675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14677 = 7'h2b == _myNewVec_14_T_3[6:0] ? myVec_43 : _GEN_14676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14678 = 7'h2c == _myNewVec_14_T_3[6:0] ? myVec_44 : _GEN_14677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14679 = 7'h2d == _myNewVec_14_T_3[6:0] ? myVec_45 : _GEN_14678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14680 = 7'h2e == _myNewVec_14_T_3[6:0] ? myVec_46 : _GEN_14679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14681 = 7'h2f == _myNewVec_14_T_3[6:0] ? myVec_47 : _GEN_14680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14682 = 7'h30 == _myNewVec_14_T_3[6:0] ? myVec_48 : _GEN_14681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14683 = 7'h31 == _myNewVec_14_T_3[6:0] ? myVec_49 : _GEN_14682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14684 = 7'h32 == _myNewVec_14_T_3[6:0] ? myVec_50 : _GEN_14683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14685 = 7'h33 == _myNewVec_14_T_3[6:0] ? myVec_51 : _GEN_14684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14686 = 7'h34 == _myNewVec_14_T_3[6:0] ? myVec_52 : _GEN_14685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14687 = 7'h35 == _myNewVec_14_T_3[6:0] ? myVec_53 : _GEN_14686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14688 = 7'h36 == _myNewVec_14_T_3[6:0] ? myVec_54 : _GEN_14687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14689 = 7'h37 == _myNewVec_14_T_3[6:0] ? myVec_55 : _GEN_14688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14690 = 7'h38 == _myNewVec_14_T_3[6:0] ? myVec_56 : _GEN_14689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14691 = 7'h39 == _myNewVec_14_T_3[6:0] ? myVec_57 : _GEN_14690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14692 = 7'h3a == _myNewVec_14_T_3[6:0] ? myVec_58 : _GEN_14691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14693 = 7'h3b == _myNewVec_14_T_3[6:0] ? myVec_59 : _GEN_14692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14694 = 7'h3c == _myNewVec_14_T_3[6:0] ? myVec_60 : _GEN_14693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14695 = 7'h3d == _myNewVec_14_T_3[6:0] ? myVec_61 : _GEN_14694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14696 = 7'h3e == _myNewVec_14_T_3[6:0] ? myVec_62 : _GEN_14695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14697 = 7'h3f == _myNewVec_14_T_3[6:0] ? myVec_63 : _GEN_14696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14698 = 7'h40 == _myNewVec_14_T_3[6:0] ? myVec_64 : _GEN_14697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14699 = 7'h41 == _myNewVec_14_T_3[6:0] ? myVec_65 : _GEN_14698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14700 = 7'h42 == _myNewVec_14_T_3[6:0] ? myVec_66 : _GEN_14699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14701 = 7'h43 == _myNewVec_14_T_3[6:0] ? myVec_67 : _GEN_14700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14702 = 7'h44 == _myNewVec_14_T_3[6:0] ? myVec_68 : _GEN_14701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14703 = 7'h45 == _myNewVec_14_T_3[6:0] ? myVec_69 : _GEN_14702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14704 = 7'h46 == _myNewVec_14_T_3[6:0] ? myVec_70 : _GEN_14703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14705 = 7'h47 == _myNewVec_14_T_3[6:0] ? myVec_71 : _GEN_14704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14706 = 7'h48 == _myNewVec_14_T_3[6:0] ? myVec_72 : _GEN_14705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14707 = 7'h49 == _myNewVec_14_T_3[6:0] ? myVec_73 : _GEN_14706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14708 = 7'h4a == _myNewVec_14_T_3[6:0] ? myVec_74 : _GEN_14707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14709 = 7'h4b == _myNewVec_14_T_3[6:0] ? myVec_75 : _GEN_14708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14710 = 7'h4c == _myNewVec_14_T_3[6:0] ? myVec_76 : _GEN_14709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14711 = 7'h4d == _myNewVec_14_T_3[6:0] ? myVec_77 : _GEN_14710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14712 = 7'h4e == _myNewVec_14_T_3[6:0] ? myVec_78 : _GEN_14711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14713 = 7'h4f == _myNewVec_14_T_3[6:0] ? myVec_79 : _GEN_14712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14714 = 7'h50 == _myNewVec_14_T_3[6:0] ? myVec_80 : _GEN_14713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14715 = 7'h51 == _myNewVec_14_T_3[6:0] ? myVec_81 : _GEN_14714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14716 = 7'h52 == _myNewVec_14_T_3[6:0] ? myVec_82 : _GEN_14715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14717 = 7'h53 == _myNewVec_14_T_3[6:0] ? myVec_83 : _GEN_14716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14718 = 7'h54 == _myNewVec_14_T_3[6:0] ? myVec_84 : _GEN_14717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14719 = 7'h55 == _myNewVec_14_T_3[6:0] ? myVec_85 : _GEN_14718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14720 = 7'h56 == _myNewVec_14_T_3[6:0] ? myVec_86 : _GEN_14719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14721 = 7'h57 == _myNewVec_14_T_3[6:0] ? myVec_87 : _GEN_14720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14722 = 7'h58 == _myNewVec_14_T_3[6:0] ? myVec_88 : _GEN_14721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14723 = 7'h59 == _myNewVec_14_T_3[6:0] ? myVec_89 : _GEN_14722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14724 = 7'h5a == _myNewVec_14_T_3[6:0] ? myVec_90 : _GEN_14723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14725 = 7'h5b == _myNewVec_14_T_3[6:0] ? myVec_91 : _GEN_14724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14726 = 7'h5c == _myNewVec_14_T_3[6:0] ? myVec_92 : _GEN_14725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14727 = 7'h5d == _myNewVec_14_T_3[6:0] ? myVec_93 : _GEN_14726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14728 = 7'h5e == _myNewVec_14_T_3[6:0] ? myVec_94 : _GEN_14727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14729 = 7'h5f == _myNewVec_14_T_3[6:0] ? myVec_95 : _GEN_14728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14730 = 7'h60 == _myNewVec_14_T_3[6:0] ? myVec_96 : _GEN_14729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14731 = 7'h61 == _myNewVec_14_T_3[6:0] ? myVec_97 : _GEN_14730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14732 = 7'h62 == _myNewVec_14_T_3[6:0] ? myVec_98 : _GEN_14731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14733 = 7'h63 == _myNewVec_14_T_3[6:0] ? myVec_99 : _GEN_14732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14734 = 7'h64 == _myNewVec_14_T_3[6:0] ? myVec_100 : _GEN_14733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14735 = 7'h65 == _myNewVec_14_T_3[6:0] ? myVec_101 : _GEN_14734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14736 = 7'h66 == _myNewVec_14_T_3[6:0] ? myVec_102 : _GEN_14735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14737 = 7'h67 == _myNewVec_14_T_3[6:0] ? myVec_103 : _GEN_14736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14738 = 7'h68 == _myNewVec_14_T_3[6:0] ? myVec_104 : _GEN_14737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14739 = 7'h69 == _myNewVec_14_T_3[6:0] ? myVec_105 : _GEN_14738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14740 = 7'h6a == _myNewVec_14_T_3[6:0] ? myVec_106 : _GEN_14739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14741 = 7'h6b == _myNewVec_14_T_3[6:0] ? myVec_107 : _GEN_14740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14742 = 7'h6c == _myNewVec_14_T_3[6:0] ? myVec_108 : _GEN_14741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14743 = 7'h6d == _myNewVec_14_T_3[6:0] ? myVec_109 : _GEN_14742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14744 = 7'h6e == _myNewVec_14_T_3[6:0] ? myVec_110 : _GEN_14743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14745 = 7'h6f == _myNewVec_14_T_3[6:0] ? myVec_111 : _GEN_14744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14746 = 7'h70 == _myNewVec_14_T_3[6:0] ? myVec_112 : _GEN_14745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14747 = 7'h71 == _myNewVec_14_T_3[6:0] ? myVec_113 : _GEN_14746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14748 = 7'h72 == _myNewVec_14_T_3[6:0] ? myVec_114 : _GEN_14747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14749 = 7'h73 == _myNewVec_14_T_3[6:0] ? myVec_115 : _GEN_14748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14750 = 7'h74 == _myNewVec_14_T_3[6:0] ? myVec_116 : _GEN_14749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14751 = 7'h75 == _myNewVec_14_T_3[6:0] ? myVec_117 : _GEN_14750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14752 = 7'h76 == _myNewVec_14_T_3[6:0] ? myVec_118 : _GEN_14751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14753 = 7'h77 == _myNewVec_14_T_3[6:0] ? myVec_119 : _GEN_14752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14754 = 7'h78 == _myNewVec_14_T_3[6:0] ? myVec_120 : _GEN_14753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14755 = 7'h79 == _myNewVec_14_T_3[6:0] ? myVec_121 : _GEN_14754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14756 = 7'h7a == _myNewVec_14_T_3[6:0] ? myVec_122 : _GEN_14755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14757 = 7'h7b == _myNewVec_14_T_3[6:0] ? myVec_123 : _GEN_14756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14758 = 7'h7c == _myNewVec_14_T_3[6:0] ? myVec_124 : _GEN_14757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14759 = 7'h7d == _myNewVec_14_T_3[6:0] ? myVec_125 : _GEN_14758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14760 = 7'h7e == _myNewVec_14_T_3[6:0] ? myVec_126 : _GEN_14759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_14 = 7'h7f == _myNewVec_14_T_3[6:0] ? myVec_127 : _GEN_14760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_13_T_3 = _myNewVec_127_T_1 + 16'h72; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_14763 = 7'h1 == _myNewVec_13_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14764 = 7'h2 == _myNewVec_13_T_3[6:0] ? myVec_2 : _GEN_14763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14765 = 7'h3 == _myNewVec_13_T_3[6:0] ? myVec_3 : _GEN_14764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14766 = 7'h4 == _myNewVec_13_T_3[6:0] ? myVec_4 : _GEN_14765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14767 = 7'h5 == _myNewVec_13_T_3[6:0] ? myVec_5 : _GEN_14766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14768 = 7'h6 == _myNewVec_13_T_3[6:0] ? myVec_6 : _GEN_14767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14769 = 7'h7 == _myNewVec_13_T_3[6:0] ? myVec_7 : _GEN_14768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14770 = 7'h8 == _myNewVec_13_T_3[6:0] ? myVec_8 : _GEN_14769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14771 = 7'h9 == _myNewVec_13_T_3[6:0] ? myVec_9 : _GEN_14770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14772 = 7'ha == _myNewVec_13_T_3[6:0] ? myVec_10 : _GEN_14771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14773 = 7'hb == _myNewVec_13_T_3[6:0] ? myVec_11 : _GEN_14772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14774 = 7'hc == _myNewVec_13_T_3[6:0] ? myVec_12 : _GEN_14773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14775 = 7'hd == _myNewVec_13_T_3[6:0] ? myVec_13 : _GEN_14774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14776 = 7'he == _myNewVec_13_T_3[6:0] ? myVec_14 : _GEN_14775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14777 = 7'hf == _myNewVec_13_T_3[6:0] ? myVec_15 : _GEN_14776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14778 = 7'h10 == _myNewVec_13_T_3[6:0] ? myVec_16 : _GEN_14777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14779 = 7'h11 == _myNewVec_13_T_3[6:0] ? myVec_17 : _GEN_14778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14780 = 7'h12 == _myNewVec_13_T_3[6:0] ? myVec_18 : _GEN_14779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14781 = 7'h13 == _myNewVec_13_T_3[6:0] ? myVec_19 : _GEN_14780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14782 = 7'h14 == _myNewVec_13_T_3[6:0] ? myVec_20 : _GEN_14781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14783 = 7'h15 == _myNewVec_13_T_3[6:0] ? myVec_21 : _GEN_14782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14784 = 7'h16 == _myNewVec_13_T_3[6:0] ? myVec_22 : _GEN_14783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14785 = 7'h17 == _myNewVec_13_T_3[6:0] ? myVec_23 : _GEN_14784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14786 = 7'h18 == _myNewVec_13_T_3[6:0] ? myVec_24 : _GEN_14785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14787 = 7'h19 == _myNewVec_13_T_3[6:0] ? myVec_25 : _GEN_14786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14788 = 7'h1a == _myNewVec_13_T_3[6:0] ? myVec_26 : _GEN_14787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14789 = 7'h1b == _myNewVec_13_T_3[6:0] ? myVec_27 : _GEN_14788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14790 = 7'h1c == _myNewVec_13_T_3[6:0] ? myVec_28 : _GEN_14789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14791 = 7'h1d == _myNewVec_13_T_3[6:0] ? myVec_29 : _GEN_14790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14792 = 7'h1e == _myNewVec_13_T_3[6:0] ? myVec_30 : _GEN_14791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14793 = 7'h1f == _myNewVec_13_T_3[6:0] ? myVec_31 : _GEN_14792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14794 = 7'h20 == _myNewVec_13_T_3[6:0] ? myVec_32 : _GEN_14793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14795 = 7'h21 == _myNewVec_13_T_3[6:0] ? myVec_33 : _GEN_14794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14796 = 7'h22 == _myNewVec_13_T_3[6:0] ? myVec_34 : _GEN_14795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14797 = 7'h23 == _myNewVec_13_T_3[6:0] ? myVec_35 : _GEN_14796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14798 = 7'h24 == _myNewVec_13_T_3[6:0] ? myVec_36 : _GEN_14797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14799 = 7'h25 == _myNewVec_13_T_3[6:0] ? myVec_37 : _GEN_14798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14800 = 7'h26 == _myNewVec_13_T_3[6:0] ? myVec_38 : _GEN_14799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14801 = 7'h27 == _myNewVec_13_T_3[6:0] ? myVec_39 : _GEN_14800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14802 = 7'h28 == _myNewVec_13_T_3[6:0] ? myVec_40 : _GEN_14801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14803 = 7'h29 == _myNewVec_13_T_3[6:0] ? myVec_41 : _GEN_14802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14804 = 7'h2a == _myNewVec_13_T_3[6:0] ? myVec_42 : _GEN_14803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14805 = 7'h2b == _myNewVec_13_T_3[6:0] ? myVec_43 : _GEN_14804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14806 = 7'h2c == _myNewVec_13_T_3[6:0] ? myVec_44 : _GEN_14805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14807 = 7'h2d == _myNewVec_13_T_3[6:0] ? myVec_45 : _GEN_14806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14808 = 7'h2e == _myNewVec_13_T_3[6:0] ? myVec_46 : _GEN_14807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14809 = 7'h2f == _myNewVec_13_T_3[6:0] ? myVec_47 : _GEN_14808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14810 = 7'h30 == _myNewVec_13_T_3[6:0] ? myVec_48 : _GEN_14809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14811 = 7'h31 == _myNewVec_13_T_3[6:0] ? myVec_49 : _GEN_14810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14812 = 7'h32 == _myNewVec_13_T_3[6:0] ? myVec_50 : _GEN_14811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14813 = 7'h33 == _myNewVec_13_T_3[6:0] ? myVec_51 : _GEN_14812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14814 = 7'h34 == _myNewVec_13_T_3[6:0] ? myVec_52 : _GEN_14813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14815 = 7'h35 == _myNewVec_13_T_3[6:0] ? myVec_53 : _GEN_14814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14816 = 7'h36 == _myNewVec_13_T_3[6:0] ? myVec_54 : _GEN_14815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14817 = 7'h37 == _myNewVec_13_T_3[6:0] ? myVec_55 : _GEN_14816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14818 = 7'h38 == _myNewVec_13_T_3[6:0] ? myVec_56 : _GEN_14817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14819 = 7'h39 == _myNewVec_13_T_3[6:0] ? myVec_57 : _GEN_14818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14820 = 7'h3a == _myNewVec_13_T_3[6:0] ? myVec_58 : _GEN_14819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14821 = 7'h3b == _myNewVec_13_T_3[6:0] ? myVec_59 : _GEN_14820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14822 = 7'h3c == _myNewVec_13_T_3[6:0] ? myVec_60 : _GEN_14821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14823 = 7'h3d == _myNewVec_13_T_3[6:0] ? myVec_61 : _GEN_14822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14824 = 7'h3e == _myNewVec_13_T_3[6:0] ? myVec_62 : _GEN_14823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14825 = 7'h3f == _myNewVec_13_T_3[6:0] ? myVec_63 : _GEN_14824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14826 = 7'h40 == _myNewVec_13_T_3[6:0] ? myVec_64 : _GEN_14825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14827 = 7'h41 == _myNewVec_13_T_3[6:0] ? myVec_65 : _GEN_14826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14828 = 7'h42 == _myNewVec_13_T_3[6:0] ? myVec_66 : _GEN_14827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14829 = 7'h43 == _myNewVec_13_T_3[6:0] ? myVec_67 : _GEN_14828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14830 = 7'h44 == _myNewVec_13_T_3[6:0] ? myVec_68 : _GEN_14829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14831 = 7'h45 == _myNewVec_13_T_3[6:0] ? myVec_69 : _GEN_14830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14832 = 7'h46 == _myNewVec_13_T_3[6:0] ? myVec_70 : _GEN_14831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14833 = 7'h47 == _myNewVec_13_T_3[6:0] ? myVec_71 : _GEN_14832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14834 = 7'h48 == _myNewVec_13_T_3[6:0] ? myVec_72 : _GEN_14833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14835 = 7'h49 == _myNewVec_13_T_3[6:0] ? myVec_73 : _GEN_14834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14836 = 7'h4a == _myNewVec_13_T_3[6:0] ? myVec_74 : _GEN_14835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14837 = 7'h4b == _myNewVec_13_T_3[6:0] ? myVec_75 : _GEN_14836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14838 = 7'h4c == _myNewVec_13_T_3[6:0] ? myVec_76 : _GEN_14837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14839 = 7'h4d == _myNewVec_13_T_3[6:0] ? myVec_77 : _GEN_14838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14840 = 7'h4e == _myNewVec_13_T_3[6:0] ? myVec_78 : _GEN_14839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14841 = 7'h4f == _myNewVec_13_T_3[6:0] ? myVec_79 : _GEN_14840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14842 = 7'h50 == _myNewVec_13_T_3[6:0] ? myVec_80 : _GEN_14841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14843 = 7'h51 == _myNewVec_13_T_3[6:0] ? myVec_81 : _GEN_14842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14844 = 7'h52 == _myNewVec_13_T_3[6:0] ? myVec_82 : _GEN_14843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14845 = 7'h53 == _myNewVec_13_T_3[6:0] ? myVec_83 : _GEN_14844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14846 = 7'h54 == _myNewVec_13_T_3[6:0] ? myVec_84 : _GEN_14845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14847 = 7'h55 == _myNewVec_13_T_3[6:0] ? myVec_85 : _GEN_14846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14848 = 7'h56 == _myNewVec_13_T_3[6:0] ? myVec_86 : _GEN_14847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14849 = 7'h57 == _myNewVec_13_T_3[6:0] ? myVec_87 : _GEN_14848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14850 = 7'h58 == _myNewVec_13_T_3[6:0] ? myVec_88 : _GEN_14849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14851 = 7'h59 == _myNewVec_13_T_3[6:0] ? myVec_89 : _GEN_14850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14852 = 7'h5a == _myNewVec_13_T_3[6:0] ? myVec_90 : _GEN_14851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14853 = 7'h5b == _myNewVec_13_T_3[6:0] ? myVec_91 : _GEN_14852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14854 = 7'h5c == _myNewVec_13_T_3[6:0] ? myVec_92 : _GEN_14853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14855 = 7'h5d == _myNewVec_13_T_3[6:0] ? myVec_93 : _GEN_14854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14856 = 7'h5e == _myNewVec_13_T_3[6:0] ? myVec_94 : _GEN_14855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14857 = 7'h5f == _myNewVec_13_T_3[6:0] ? myVec_95 : _GEN_14856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14858 = 7'h60 == _myNewVec_13_T_3[6:0] ? myVec_96 : _GEN_14857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14859 = 7'h61 == _myNewVec_13_T_3[6:0] ? myVec_97 : _GEN_14858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14860 = 7'h62 == _myNewVec_13_T_3[6:0] ? myVec_98 : _GEN_14859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14861 = 7'h63 == _myNewVec_13_T_3[6:0] ? myVec_99 : _GEN_14860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14862 = 7'h64 == _myNewVec_13_T_3[6:0] ? myVec_100 : _GEN_14861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14863 = 7'h65 == _myNewVec_13_T_3[6:0] ? myVec_101 : _GEN_14862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14864 = 7'h66 == _myNewVec_13_T_3[6:0] ? myVec_102 : _GEN_14863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14865 = 7'h67 == _myNewVec_13_T_3[6:0] ? myVec_103 : _GEN_14864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14866 = 7'h68 == _myNewVec_13_T_3[6:0] ? myVec_104 : _GEN_14865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14867 = 7'h69 == _myNewVec_13_T_3[6:0] ? myVec_105 : _GEN_14866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14868 = 7'h6a == _myNewVec_13_T_3[6:0] ? myVec_106 : _GEN_14867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14869 = 7'h6b == _myNewVec_13_T_3[6:0] ? myVec_107 : _GEN_14868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14870 = 7'h6c == _myNewVec_13_T_3[6:0] ? myVec_108 : _GEN_14869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14871 = 7'h6d == _myNewVec_13_T_3[6:0] ? myVec_109 : _GEN_14870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14872 = 7'h6e == _myNewVec_13_T_3[6:0] ? myVec_110 : _GEN_14871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14873 = 7'h6f == _myNewVec_13_T_3[6:0] ? myVec_111 : _GEN_14872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14874 = 7'h70 == _myNewVec_13_T_3[6:0] ? myVec_112 : _GEN_14873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14875 = 7'h71 == _myNewVec_13_T_3[6:0] ? myVec_113 : _GEN_14874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14876 = 7'h72 == _myNewVec_13_T_3[6:0] ? myVec_114 : _GEN_14875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14877 = 7'h73 == _myNewVec_13_T_3[6:0] ? myVec_115 : _GEN_14876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14878 = 7'h74 == _myNewVec_13_T_3[6:0] ? myVec_116 : _GEN_14877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14879 = 7'h75 == _myNewVec_13_T_3[6:0] ? myVec_117 : _GEN_14878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14880 = 7'h76 == _myNewVec_13_T_3[6:0] ? myVec_118 : _GEN_14879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14881 = 7'h77 == _myNewVec_13_T_3[6:0] ? myVec_119 : _GEN_14880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14882 = 7'h78 == _myNewVec_13_T_3[6:0] ? myVec_120 : _GEN_14881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14883 = 7'h79 == _myNewVec_13_T_3[6:0] ? myVec_121 : _GEN_14882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14884 = 7'h7a == _myNewVec_13_T_3[6:0] ? myVec_122 : _GEN_14883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14885 = 7'h7b == _myNewVec_13_T_3[6:0] ? myVec_123 : _GEN_14884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14886 = 7'h7c == _myNewVec_13_T_3[6:0] ? myVec_124 : _GEN_14885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14887 = 7'h7d == _myNewVec_13_T_3[6:0] ? myVec_125 : _GEN_14886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14888 = 7'h7e == _myNewVec_13_T_3[6:0] ? myVec_126 : _GEN_14887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_13 = 7'h7f == _myNewVec_13_T_3[6:0] ? myVec_127 : _GEN_14888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_12_T_3 = _myNewVec_127_T_1 + 16'h73; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_14891 = 7'h1 == _myNewVec_12_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14892 = 7'h2 == _myNewVec_12_T_3[6:0] ? myVec_2 : _GEN_14891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14893 = 7'h3 == _myNewVec_12_T_3[6:0] ? myVec_3 : _GEN_14892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14894 = 7'h4 == _myNewVec_12_T_3[6:0] ? myVec_4 : _GEN_14893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14895 = 7'h5 == _myNewVec_12_T_3[6:0] ? myVec_5 : _GEN_14894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14896 = 7'h6 == _myNewVec_12_T_3[6:0] ? myVec_6 : _GEN_14895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14897 = 7'h7 == _myNewVec_12_T_3[6:0] ? myVec_7 : _GEN_14896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14898 = 7'h8 == _myNewVec_12_T_3[6:0] ? myVec_8 : _GEN_14897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14899 = 7'h9 == _myNewVec_12_T_3[6:0] ? myVec_9 : _GEN_14898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14900 = 7'ha == _myNewVec_12_T_3[6:0] ? myVec_10 : _GEN_14899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14901 = 7'hb == _myNewVec_12_T_3[6:0] ? myVec_11 : _GEN_14900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14902 = 7'hc == _myNewVec_12_T_3[6:0] ? myVec_12 : _GEN_14901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14903 = 7'hd == _myNewVec_12_T_3[6:0] ? myVec_13 : _GEN_14902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14904 = 7'he == _myNewVec_12_T_3[6:0] ? myVec_14 : _GEN_14903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14905 = 7'hf == _myNewVec_12_T_3[6:0] ? myVec_15 : _GEN_14904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14906 = 7'h10 == _myNewVec_12_T_3[6:0] ? myVec_16 : _GEN_14905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14907 = 7'h11 == _myNewVec_12_T_3[6:0] ? myVec_17 : _GEN_14906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14908 = 7'h12 == _myNewVec_12_T_3[6:0] ? myVec_18 : _GEN_14907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14909 = 7'h13 == _myNewVec_12_T_3[6:0] ? myVec_19 : _GEN_14908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14910 = 7'h14 == _myNewVec_12_T_3[6:0] ? myVec_20 : _GEN_14909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14911 = 7'h15 == _myNewVec_12_T_3[6:0] ? myVec_21 : _GEN_14910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14912 = 7'h16 == _myNewVec_12_T_3[6:0] ? myVec_22 : _GEN_14911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14913 = 7'h17 == _myNewVec_12_T_3[6:0] ? myVec_23 : _GEN_14912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14914 = 7'h18 == _myNewVec_12_T_3[6:0] ? myVec_24 : _GEN_14913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14915 = 7'h19 == _myNewVec_12_T_3[6:0] ? myVec_25 : _GEN_14914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14916 = 7'h1a == _myNewVec_12_T_3[6:0] ? myVec_26 : _GEN_14915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14917 = 7'h1b == _myNewVec_12_T_3[6:0] ? myVec_27 : _GEN_14916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14918 = 7'h1c == _myNewVec_12_T_3[6:0] ? myVec_28 : _GEN_14917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14919 = 7'h1d == _myNewVec_12_T_3[6:0] ? myVec_29 : _GEN_14918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14920 = 7'h1e == _myNewVec_12_T_3[6:0] ? myVec_30 : _GEN_14919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14921 = 7'h1f == _myNewVec_12_T_3[6:0] ? myVec_31 : _GEN_14920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14922 = 7'h20 == _myNewVec_12_T_3[6:0] ? myVec_32 : _GEN_14921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14923 = 7'h21 == _myNewVec_12_T_3[6:0] ? myVec_33 : _GEN_14922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14924 = 7'h22 == _myNewVec_12_T_3[6:0] ? myVec_34 : _GEN_14923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14925 = 7'h23 == _myNewVec_12_T_3[6:0] ? myVec_35 : _GEN_14924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14926 = 7'h24 == _myNewVec_12_T_3[6:0] ? myVec_36 : _GEN_14925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14927 = 7'h25 == _myNewVec_12_T_3[6:0] ? myVec_37 : _GEN_14926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14928 = 7'h26 == _myNewVec_12_T_3[6:0] ? myVec_38 : _GEN_14927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14929 = 7'h27 == _myNewVec_12_T_3[6:0] ? myVec_39 : _GEN_14928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14930 = 7'h28 == _myNewVec_12_T_3[6:0] ? myVec_40 : _GEN_14929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14931 = 7'h29 == _myNewVec_12_T_3[6:0] ? myVec_41 : _GEN_14930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14932 = 7'h2a == _myNewVec_12_T_3[6:0] ? myVec_42 : _GEN_14931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14933 = 7'h2b == _myNewVec_12_T_3[6:0] ? myVec_43 : _GEN_14932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14934 = 7'h2c == _myNewVec_12_T_3[6:0] ? myVec_44 : _GEN_14933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14935 = 7'h2d == _myNewVec_12_T_3[6:0] ? myVec_45 : _GEN_14934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14936 = 7'h2e == _myNewVec_12_T_3[6:0] ? myVec_46 : _GEN_14935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14937 = 7'h2f == _myNewVec_12_T_3[6:0] ? myVec_47 : _GEN_14936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14938 = 7'h30 == _myNewVec_12_T_3[6:0] ? myVec_48 : _GEN_14937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14939 = 7'h31 == _myNewVec_12_T_3[6:0] ? myVec_49 : _GEN_14938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14940 = 7'h32 == _myNewVec_12_T_3[6:0] ? myVec_50 : _GEN_14939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14941 = 7'h33 == _myNewVec_12_T_3[6:0] ? myVec_51 : _GEN_14940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14942 = 7'h34 == _myNewVec_12_T_3[6:0] ? myVec_52 : _GEN_14941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14943 = 7'h35 == _myNewVec_12_T_3[6:0] ? myVec_53 : _GEN_14942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14944 = 7'h36 == _myNewVec_12_T_3[6:0] ? myVec_54 : _GEN_14943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14945 = 7'h37 == _myNewVec_12_T_3[6:0] ? myVec_55 : _GEN_14944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14946 = 7'h38 == _myNewVec_12_T_3[6:0] ? myVec_56 : _GEN_14945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14947 = 7'h39 == _myNewVec_12_T_3[6:0] ? myVec_57 : _GEN_14946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14948 = 7'h3a == _myNewVec_12_T_3[6:0] ? myVec_58 : _GEN_14947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14949 = 7'h3b == _myNewVec_12_T_3[6:0] ? myVec_59 : _GEN_14948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14950 = 7'h3c == _myNewVec_12_T_3[6:0] ? myVec_60 : _GEN_14949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14951 = 7'h3d == _myNewVec_12_T_3[6:0] ? myVec_61 : _GEN_14950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14952 = 7'h3e == _myNewVec_12_T_3[6:0] ? myVec_62 : _GEN_14951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14953 = 7'h3f == _myNewVec_12_T_3[6:0] ? myVec_63 : _GEN_14952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14954 = 7'h40 == _myNewVec_12_T_3[6:0] ? myVec_64 : _GEN_14953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14955 = 7'h41 == _myNewVec_12_T_3[6:0] ? myVec_65 : _GEN_14954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14956 = 7'h42 == _myNewVec_12_T_3[6:0] ? myVec_66 : _GEN_14955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14957 = 7'h43 == _myNewVec_12_T_3[6:0] ? myVec_67 : _GEN_14956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14958 = 7'h44 == _myNewVec_12_T_3[6:0] ? myVec_68 : _GEN_14957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14959 = 7'h45 == _myNewVec_12_T_3[6:0] ? myVec_69 : _GEN_14958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14960 = 7'h46 == _myNewVec_12_T_3[6:0] ? myVec_70 : _GEN_14959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14961 = 7'h47 == _myNewVec_12_T_3[6:0] ? myVec_71 : _GEN_14960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14962 = 7'h48 == _myNewVec_12_T_3[6:0] ? myVec_72 : _GEN_14961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14963 = 7'h49 == _myNewVec_12_T_3[6:0] ? myVec_73 : _GEN_14962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14964 = 7'h4a == _myNewVec_12_T_3[6:0] ? myVec_74 : _GEN_14963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14965 = 7'h4b == _myNewVec_12_T_3[6:0] ? myVec_75 : _GEN_14964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14966 = 7'h4c == _myNewVec_12_T_3[6:0] ? myVec_76 : _GEN_14965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14967 = 7'h4d == _myNewVec_12_T_3[6:0] ? myVec_77 : _GEN_14966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14968 = 7'h4e == _myNewVec_12_T_3[6:0] ? myVec_78 : _GEN_14967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14969 = 7'h4f == _myNewVec_12_T_3[6:0] ? myVec_79 : _GEN_14968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14970 = 7'h50 == _myNewVec_12_T_3[6:0] ? myVec_80 : _GEN_14969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14971 = 7'h51 == _myNewVec_12_T_3[6:0] ? myVec_81 : _GEN_14970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14972 = 7'h52 == _myNewVec_12_T_3[6:0] ? myVec_82 : _GEN_14971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14973 = 7'h53 == _myNewVec_12_T_3[6:0] ? myVec_83 : _GEN_14972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14974 = 7'h54 == _myNewVec_12_T_3[6:0] ? myVec_84 : _GEN_14973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14975 = 7'h55 == _myNewVec_12_T_3[6:0] ? myVec_85 : _GEN_14974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14976 = 7'h56 == _myNewVec_12_T_3[6:0] ? myVec_86 : _GEN_14975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14977 = 7'h57 == _myNewVec_12_T_3[6:0] ? myVec_87 : _GEN_14976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14978 = 7'h58 == _myNewVec_12_T_3[6:0] ? myVec_88 : _GEN_14977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14979 = 7'h59 == _myNewVec_12_T_3[6:0] ? myVec_89 : _GEN_14978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14980 = 7'h5a == _myNewVec_12_T_3[6:0] ? myVec_90 : _GEN_14979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14981 = 7'h5b == _myNewVec_12_T_3[6:0] ? myVec_91 : _GEN_14980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14982 = 7'h5c == _myNewVec_12_T_3[6:0] ? myVec_92 : _GEN_14981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14983 = 7'h5d == _myNewVec_12_T_3[6:0] ? myVec_93 : _GEN_14982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14984 = 7'h5e == _myNewVec_12_T_3[6:0] ? myVec_94 : _GEN_14983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14985 = 7'h5f == _myNewVec_12_T_3[6:0] ? myVec_95 : _GEN_14984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14986 = 7'h60 == _myNewVec_12_T_3[6:0] ? myVec_96 : _GEN_14985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14987 = 7'h61 == _myNewVec_12_T_3[6:0] ? myVec_97 : _GEN_14986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14988 = 7'h62 == _myNewVec_12_T_3[6:0] ? myVec_98 : _GEN_14987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14989 = 7'h63 == _myNewVec_12_T_3[6:0] ? myVec_99 : _GEN_14988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14990 = 7'h64 == _myNewVec_12_T_3[6:0] ? myVec_100 : _GEN_14989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14991 = 7'h65 == _myNewVec_12_T_3[6:0] ? myVec_101 : _GEN_14990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14992 = 7'h66 == _myNewVec_12_T_3[6:0] ? myVec_102 : _GEN_14991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14993 = 7'h67 == _myNewVec_12_T_3[6:0] ? myVec_103 : _GEN_14992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14994 = 7'h68 == _myNewVec_12_T_3[6:0] ? myVec_104 : _GEN_14993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14995 = 7'h69 == _myNewVec_12_T_3[6:0] ? myVec_105 : _GEN_14994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14996 = 7'h6a == _myNewVec_12_T_3[6:0] ? myVec_106 : _GEN_14995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14997 = 7'h6b == _myNewVec_12_T_3[6:0] ? myVec_107 : _GEN_14996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14998 = 7'h6c == _myNewVec_12_T_3[6:0] ? myVec_108 : _GEN_14997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_14999 = 7'h6d == _myNewVec_12_T_3[6:0] ? myVec_109 : _GEN_14998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15000 = 7'h6e == _myNewVec_12_T_3[6:0] ? myVec_110 : _GEN_14999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15001 = 7'h6f == _myNewVec_12_T_3[6:0] ? myVec_111 : _GEN_15000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15002 = 7'h70 == _myNewVec_12_T_3[6:0] ? myVec_112 : _GEN_15001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15003 = 7'h71 == _myNewVec_12_T_3[6:0] ? myVec_113 : _GEN_15002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15004 = 7'h72 == _myNewVec_12_T_3[6:0] ? myVec_114 : _GEN_15003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15005 = 7'h73 == _myNewVec_12_T_3[6:0] ? myVec_115 : _GEN_15004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15006 = 7'h74 == _myNewVec_12_T_3[6:0] ? myVec_116 : _GEN_15005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15007 = 7'h75 == _myNewVec_12_T_3[6:0] ? myVec_117 : _GEN_15006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15008 = 7'h76 == _myNewVec_12_T_3[6:0] ? myVec_118 : _GEN_15007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15009 = 7'h77 == _myNewVec_12_T_3[6:0] ? myVec_119 : _GEN_15008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15010 = 7'h78 == _myNewVec_12_T_3[6:0] ? myVec_120 : _GEN_15009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15011 = 7'h79 == _myNewVec_12_T_3[6:0] ? myVec_121 : _GEN_15010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15012 = 7'h7a == _myNewVec_12_T_3[6:0] ? myVec_122 : _GEN_15011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15013 = 7'h7b == _myNewVec_12_T_3[6:0] ? myVec_123 : _GEN_15012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15014 = 7'h7c == _myNewVec_12_T_3[6:0] ? myVec_124 : _GEN_15013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15015 = 7'h7d == _myNewVec_12_T_3[6:0] ? myVec_125 : _GEN_15014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15016 = 7'h7e == _myNewVec_12_T_3[6:0] ? myVec_126 : _GEN_15015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_12 = 7'h7f == _myNewVec_12_T_3[6:0] ? myVec_127 : _GEN_15016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_11_T_3 = _myNewVec_127_T_1 + 16'h74; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_15019 = 7'h1 == _myNewVec_11_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15020 = 7'h2 == _myNewVec_11_T_3[6:0] ? myVec_2 : _GEN_15019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15021 = 7'h3 == _myNewVec_11_T_3[6:0] ? myVec_3 : _GEN_15020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15022 = 7'h4 == _myNewVec_11_T_3[6:0] ? myVec_4 : _GEN_15021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15023 = 7'h5 == _myNewVec_11_T_3[6:0] ? myVec_5 : _GEN_15022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15024 = 7'h6 == _myNewVec_11_T_3[6:0] ? myVec_6 : _GEN_15023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15025 = 7'h7 == _myNewVec_11_T_3[6:0] ? myVec_7 : _GEN_15024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15026 = 7'h8 == _myNewVec_11_T_3[6:0] ? myVec_8 : _GEN_15025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15027 = 7'h9 == _myNewVec_11_T_3[6:0] ? myVec_9 : _GEN_15026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15028 = 7'ha == _myNewVec_11_T_3[6:0] ? myVec_10 : _GEN_15027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15029 = 7'hb == _myNewVec_11_T_3[6:0] ? myVec_11 : _GEN_15028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15030 = 7'hc == _myNewVec_11_T_3[6:0] ? myVec_12 : _GEN_15029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15031 = 7'hd == _myNewVec_11_T_3[6:0] ? myVec_13 : _GEN_15030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15032 = 7'he == _myNewVec_11_T_3[6:0] ? myVec_14 : _GEN_15031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15033 = 7'hf == _myNewVec_11_T_3[6:0] ? myVec_15 : _GEN_15032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15034 = 7'h10 == _myNewVec_11_T_3[6:0] ? myVec_16 : _GEN_15033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15035 = 7'h11 == _myNewVec_11_T_3[6:0] ? myVec_17 : _GEN_15034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15036 = 7'h12 == _myNewVec_11_T_3[6:0] ? myVec_18 : _GEN_15035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15037 = 7'h13 == _myNewVec_11_T_3[6:0] ? myVec_19 : _GEN_15036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15038 = 7'h14 == _myNewVec_11_T_3[6:0] ? myVec_20 : _GEN_15037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15039 = 7'h15 == _myNewVec_11_T_3[6:0] ? myVec_21 : _GEN_15038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15040 = 7'h16 == _myNewVec_11_T_3[6:0] ? myVec_22 : _GEN_15039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15041 = 7'h17 == _myNewVec_11_T_3[6:0] ? myVec_23 : _GEN_15040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15042 = 7'h18 == _myNewVec_11_T_3[6:0] ? myVec_24 : _GEN_15041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15043 = 7'h19 == _myNewVec_11_T_3[6:0] ? myVec_25 : _GEN_15042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15044 = 7'h1a == _myNewVec_11_T_3[6:0] ? myVec_26 : _GEN_15043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15045 = 7'h1b == _myNewVec_11_T_3[6:0] ? myVec_27 : _GEN_15044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15046 = 7'h1c == _myNewVec_11_T_3[6:0] ? myVec_28 : _GEN_15045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15047 = 7'h1d == _myNewVec_11_T_3[6:0] ? myVec_29 : _GEN_15046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15048 = 7'h1e == _myNewVec_11_T_3[6:0] ? myVec_30 : _GEN_15047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15049 = 7'h1f == _myNewVec_11_T_3[6:0] ? myVec_31 : _GEN_15048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15050 = 7'h20 == _myNewVec_11_T_3[6:0] ? myVec_32 : _GEN_15049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15051 = 7'h21 == _myNewVec_11_T_3[6:0] ? myVec_33 : _GEN_15050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15052 = 7'h22 == _myNewVec_11_T_3[6:0] ? myVec_34 : _GEN_15051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15053 = 7'h23 == _myNewVec_11_T_3[6:0] ? myVec_35 : _GEN_15052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15054 = 7'h24 == _myNewVec_11_T_3[6:0] ? myVec_36 : _GEN_15053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15055 = 7'h25 == _myNewVec_11_T_3[6:0] ? myVec_37 : _GEN_15054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15056 = 7'h26 == _myNewVec_11_T_3[6:0] ? myVec_38 : _GEN_15055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15057 = 7'h27 == _myNewVec_11_T_3[6:0] ? myVec_39 : _GEN_15056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15058 = 7'h28 == _myNewVec_11_T_3[6:0] ? myVec_40 : _GEN_15057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15059 = 7'h29 == _myNewVec_11_T_3[6:0] ? myVec_41 : _GEN_15058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15060 = 7'h2a == _myNewVec_11_T_3[6:0] ? myVec_42 : _GEN_15059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15061 = 7'h2b == _myNewVec_11_T_3[6:0] ? myVec_43 : _GEN_15060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15062 = 7'h2c == _myNewVec_11_T_3[6:0] ? myVec_44 : _GEN_15061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15063 = 7'h2d == _myNewVec_11_T_3[6:0] ? myVec_45 : _GEN_15062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15064 = 7'h2e == _myNewVec_11_T_3[6:0] ? myVec_46 : _GEN_15063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15065 = 7'h2f == _myNewVec_11_T_3[6:0] ? myVec_47 : _GEN_15064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15066 = 7'h30 == _myNewVec_11_T_3[6:0] ? myVec_48 : _GEN_15065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15067 = 7'h31 == _myNewVec_11_T_3[6:0] ? myVec_49 : _GEN_15066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15068 = 7'h32 == _myNewVec_11_T_3[6:0] ? myVec_50 : _GEN_15067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15069 = 7'h33 == _myNewVec_11_T_3[6:0] ? myVec_51 : _GEN_15068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15070 = 7'h34 == _myNewVec_11_T_3[6:0] ? myVec_52 : _GEN_15069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15071 = 7'h35 == _myNewVec_11_T_3[6:0] ? myVec_53 : _GEN_15070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15072 = 7'h36 == _myNewVec_11_T_3[6:0] ? myVec_54 : _GEN_15071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15073 = 7'h37 == _myNewVec_11_T_3[6:0] ? myVec_55 : _GEN_15072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15074 = 7'h38 == _myNewVec_11_T_3[6:0] ? myVec_56 : _GEN_15073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15075 = 7'h39 == _myNewVec_11_T_3[6:0] ? myVec_57 : _GEN_15074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15076 = 7'h3a == _myNewVec_11_T_3[6:0] ? myVec_58 : _GEN_15075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15077 = 7'h3b == _myNewVec_11_T_3[6:0] ? myVec_59 : _GEN_15076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15078 = 7'h3c == _myNewVec_11_T_3[6:0] ? myVec_60 : _GEN_15077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15079 = 7'h3d == _myNewVec_11_T_3[6:0] ? myVec_61 : _GEN_15078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15080 = 7'h3e == _myNewVec_11_T_3[6:0] ? myVec_62 : _GEN_15079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15081 = 7'h3f == _myNewVec_11_T_3[6:0] ? myVec_63 : _GEN_15080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15082 = 7'h40 == _myNewVec_11_T_3[6:0] ? myVec_64 : _GEN_15081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15083 = 7'h41 == _myNewVec_11_T_3[6:0] ? myVec_65 : _GEN_15082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15084 = 7'h42 == _myNewVec_11_T_3[6:0] ? myVec_66 : _GEN_15083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15085 = 7'h43 == _myNewVec_11_T_3[6:0] ? myVec_67 : _GEN_15084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15086 = 7'h44 == _myNewVec_11_T_3[6:0] ? myVec_68 : _GEN_15085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15087 = 7'h45 == _myNewVec_11_T_3[6:0] ? myVec_69 : _GEN_15086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15088 = 7'h46 == _myNewVec_11_T_3[6:0] ? myVec_70 : _GEN_15087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15089 = 7'h47 == _myNewVec_11_T_3[6:0] ? myVec_71 : _GEN_15088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15090 = 7'h48 == _myNewVec_11_T_3[6:0] ? myVec_72 : _GEN_15089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15091 = 7'h49 == _myNewVec_11_T_3[6:0] ? myVec_73 : _GEN_15090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15092 = 7'h4a == _myNewVec_11_T_3[6:0] ? myVec_74 : _GEN_15091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15093 = 7'h4b == _myNewVec_11_T_3[6:0] ? myVec_75 : _GEN_15092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15094 = 7'h4c == _myNewVec_11_T_3[6:0] ? myVec_76 : _GEN_15093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15095 = 7'h4d == _myNewVec_11_T_3[6:0] ? myVec_77 : _GEN_15094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15096 = 7'h4e == _myNewVec_11_T_3[6:0] ? myVec_78 : _GEN_15095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15097 = 7'h4f == _myNewVec_11_T_3[6:0] ? myVec_79 : _GEN_15096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15098 = 7'h50 == _myNewVec_11_T_3[6:0] ? myVec_80 : _GEN_15097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15099 = 7'h51 == _myNewVec_11_T_3[6:0] ? myVec_81 : _GEN_15098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15100 = 7'h52 == _myNewVec_11_T_3[6:0] ? myVec_82 : _GEN_15099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15101 = 7'h53 == _myNewVec_11_T_3[6:0] ? myVec_83 : _GEN_15100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15102 = 7'h54 == _myNewVec_11_T_3[6:0] ? myVec_84 : _GEN_15101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15103 = 7'h55 == _myNewVec_11_T_3[6:0] ? myVec_85 : _GEN_15102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15104 = 7'h56 == _myNewVec_11_T_3[6:0] ? myVec_86 : _GEN_15103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15105 = 7'h57 == _myNewVec_11_T_3[6:0] ? myVec_87 : _GEN_15104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15106 = 7'h58 == _myNewVec_11_T_3[6:0] ? myVec_88 : _GEN_15105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15107 = 7'h59 == _myNewVec_11_T_3[6:0] ? myVec_89 : _GEN_15106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15108 = 7'h5a == _myNewVec_11_T_3[6:0] ? myVec_90 : _GEN_15107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15109 = 7'h5b == _myNewVec_11_T_3[6:0] ? myVec_91 : _GEN_15108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15110 = 7'h5c == _myNewVec_11_T_3[6:0] ? myVec_92 : _GEN_15109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15111 = 7'h5d == _myNewVec_11_T_3[6:0] ? myVec_93 : _GEN_15110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15112 = 7'h5e == _myNewVec_11_T_3[6:0] ? myVec_94 : _GEN_15111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15113 = 7'h5f == _myNewVec_11_T_3[6:0] ? myVec_95 : _GEN_15112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15114 = 7'h60 == _myNewVec_11_T_3[6:0] ? myVec_96 : _GEN_15113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15115 = 7'h61 == _myNewVec_11_T_3[6:0] ? myVec_97 : _GEN_15114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15116 = 7'h62 == _myNewVec_11_T_3[6:0] ? myVec_98 : _GEN_15115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15117 = 7'h63 == _myNewVec_11_T_3[6:0] ? myVec_99 : _GEN_15116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15118 = 7'h64 == _myNewVec_11_T_3[6:0] ? myVec_100 : _GEN_15117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15119 = 7'h65 == _myNewVec_11_T_3[6:0] ? myVec_101 : _GEN_15118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15120 = 7'h66 == _myNewVec_11_T_3[6:0] ? myVec_102 : _GEN_15119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15121 = 7'h67 == _myNewVec_11_T_3[6:0] ? myVec_103 : _GEN_15120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15122 = 7'h68 == _myNewVec_11_T_3[6:0] ? myVec_104 : _GEN_15121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15123 = 7'h69 == _myNewVec_11_T_3[6:0] ? myVec_105 : _GEN_15122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15124 = 7'h6a == _myNewVec_11_T_3[6:0] ? myVec_106 : _GEN_15123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15125 = 7'h6b == _myNewVec_11_T_3[6:0] ? myVec_107 : _GEN_15124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15126 = 7'h6c == _myNewVec_11_T_3[6:0] ? myVec_108 : _GEN_15125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15127 = 7'h6d == _myNewVec_11_T_3[6:0] ? myVec_109 : _GEN_15126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15128 = 7'h6e == _myNewVec_11_T_3[6:0] ? myVec_110 : _GEN_15127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15129 = 7'h6f == _myNewVec_11_T_3[6:0] ? myVec_111 : _GEN_15128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15130 = 7'h70 == _myNewVec_11_T_3[6:0] ? myVec_112 : _GEN_15129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15131 = 7'h71 == _myNewVec_11_T_3[6:0] ? myVec_113 : _GEN_15130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15132 = 7'h72 == _myNewVec_11_T_3[6:0] ? myVec_114 : _GEN_15131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15133 = 7'h73 == _myNewVec_11_T_3[6:0] ? myVec_115 : _GEN_15132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15134 = 7'h74 == _myNewVec_11_T_3[6:0] ? myVec_116 : _GEN_15133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15135 = 7'h75 == _myNewVec_11_T_3[6:0] ? myVec_117 : _GEN_15134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15136 = 7'h76 == _myNewVec_11_T_3[6:0] ? myVec_118 : _GEN_15135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15137 = 7'h77 == _myNewVec_11_T_3[6:0] ? myVec_119 : _GEN_15136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15138 = 7'h78 == _myNewVec_11_T_3[6:0] ? myVec_120 : _GEN_15137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15139 = 7'h79 == _myNewVec_11_T_3[6:0] ? myVec_121 : _GEN_15138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15140 = 7'h7a == _myNewVec_11_T_3[6:0] ? myVec_122 : _GEN_15139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15141 = 7'h7b == _myNewVec_11_T_3[6:0] ? myVec_123 : _GEN_15140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15142 = 7'h7c == _myNewVec_11_T_3[6:0] ? myVec_124 : _GEN_15141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15143 = 7'h7d == _myNewVec_11_T_3[6:0] ? myVec_125 : _GEN_15142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15144 = 7'h7e == _myNewVec_11_T_3[6:0] ? myVec_126 : _GEN_15143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_11 = 7'h7f == _myNewVec_11_T_3[6:0] ? myVec_127 : _GEN_15144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_10_T_3 = _myNewVec_127_T_1 + 16'h75; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_15147 = 7'h1 == _myNewVec_10_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15148 = 7'h2 == _myNewVec_10_T_3[6:0] ? myVec_2 : _GEN_15147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15149 = 7'h3 == _myNewVec_10_T_3[6:0] ? myVec_3 : _GEN_15148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15150 = 7'h4 == _myNewVec_10_T_3[6:0] ? myVec_4 : _GEN_15149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15151 = 7'h5 == _myNewVec_10_T_3[6:0] ? myVec_5 : _GEN_15150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15152 = 7'h6 == _myNewVec_10_T_3[6:0] ? myVec_6 : _GEN_15151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15153 = 7'h7 == _myNewVec_10_T_3[6:0] ? myVec_7 : _GEN_15152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15154 = 7'h8 == _myNewVec_10_T_3[6:0] ? myVec_8 : _GEN_15153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15155 = 7'h9 == _myNewVec_10_T_3[6:0] ? myVec_9 : _GEN_15154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15156 = 7'ha == _myNewVec_10_T_3[6:0] ? myVec_10 : _GEN_15155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15157 = 7'hb == _myNewVec_10_T_3[6:0] ? myVec_11 : _GEN_15156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15158 = 7'hc == _myNewVec_10_T_3[6:0] ? myVec_12 : _GEN_15157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15159 = 7'hd == _myNewVec_10_T_3[6:0] ? myVec_13 : _GEN_15158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15160 = 7'he == _myNewVec_10_T_3[6:0] ? myVec_14 : _GEN_15159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15161 = 7'hf == _myNewVec_10_T_3[6:0] ? myVec_15 : _GEN_15160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15162 = 7'h10 == _myNewVec_10_T_3[6:0] ? myVec_16 : _GEN_15161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15163 = 7'h11 == _myNewVec_10_T_3[6:0] ? myVec_17 : _GEN_15162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15164 = 7'h12 == _myNewVec_10_T_3[6:0] ? myVec_18 : _GEN_15163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15165 = 7'h13 == _myNewVec_10_T_3[6:0] ? myVec_19 : _GEN_15164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15166 = 7'h14 == _myNewVec_10_T_3[6:0] ? myVec_20 : _GEN_15165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15167 = 7'h15 == _myNewVec_10_T_3[6:0] ? myVec_21 : _GEN_15166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15168 = 7'h16 == _myNewVec_10_T_3[6:0] ? myVec_22 : _GEN_15167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15169 = 7'h17 == _myNewVec_10_T_3[6:0] ? myVec_23 : _GEN_15168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15170 = 7'h18 == _myNewVec_10_T_3[6:0] ? myVec_24 : _GEN_15169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15171 = 7'h19 == _myNewVec_10_T_3[6:0] ? myVec_25 : _GEN_15170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15172 = 7'h1a == _myNewVec_10_T_3[6:0] ? myVec_26 : _GEN_15171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15173 = 7'h1b == _myNewVec_10_T_3[6:0] ? myVec_27 : _GEN_15172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15174 = 7'h1c == _myNewVec_10_T_3[6:0] ? myVec_28 : _GEN_15173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15175 = 7'h1d == _myNewVec_10_T_3[6:0] ? myVec_29 : _GEN_15174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15176 = 7'h1e == _myNewVec_10_T_3[6:0] ? myVec_30 : _GEN_15175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15177 = 7'h1f == _myNewVec_10_T_3[6:0] ? myVec_31 : _GEN_15176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15178 = 7'h20 == _myNewVec_10_T_3[6:0] ? myVec_32 : _GEN_15177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15179 = 7'h21 == _myNewVec_10_T_3[6:0] ? myVec_33 : _GEN_15178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15180 = 7'h22 == _myNewVec_10_T_3[6:0] ? myVec_34 : _GEN_15179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15181 = 7'h23 == _myNewVec_10_T_3[6:0] ? myVec_35 : _GEN_15180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15182 = 7'h24 == _myNewVec_10_T_3[6:0] ? myVec_36 : _GEN_15181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15183 = 7'h25 == _myNewVec_10_T_3[6:0] ? myVec_37 : _GEN_15182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15184 = 7'h26 == _myNewVec_10_T_3[6:0] ? myVec_38 : _GEN_15183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15185 = 7'h27 == _myNewVec_10_T_3[6:0] ? myVec_39 : _GEN_15184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15186 = 7'h28 == _myNewVec_10_T_3[6:0] ? myVec_40 : _GEN_15185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15187 = 7'h29 == _myNewVec_10_T_3[6:0] ? myVec_41 : _GEN_15186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15188 = 7'h2a == _myNewVec_10_T_3[6:0] ? myVec_42 : _GEN_15187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15189 = 7'h2b == _myNewVec_10_T_3[6:0] ? myVec_43 : _GEN_15188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15190 = 7'h2c == _myNewVec_10_T_3[6:0] ? myVec_44 : _GEN_15189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15191 = 7'h2d == _myNewVec_10_T_3[6:0] ? myVec_45 : _GEN_15190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15192 = 7'h2e == _myNewVec_10_T_3[6:0] ? myVec_46 : _GEN_15191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15193 = 7'h2f == _myNewVec_10_T_3[6:0] ? myVec_47 : _GEN_15192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15194 = 7'h30 == _myNewVec_10_T_3[6:0] ? myVec_48 : _GEN_15193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15195 = 7'h31 == _myNewVec_10_T_3[6:0] ? myVec_49 : _GEN_15194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15196 = 7'h32 == _myNewVec_10_T_3[6:0] ? myVec_50 : _GEN_15195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15197 = 7'h33 == _myNewVec_10_T_3[6:0] ? myVec_51 : _GEN_15196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15198 = 7'h34 == _myNewVec_10_T_3[6:0] ? myVec_52 : _GEN_15197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15199 = 7'h35 == _myNewVec_10_T_3[6:0] ? myVec_53 : _GEN_15198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15200 = 7'h36 == _myNewVec_10_T_3[6:0] ? myVec_54 : _GEN_15199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15201 = 7'h37 == _myNewVec_10_T_3[6:0] ? myVec_55 : _GEN_15200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15202 = 7'h38 == _myNewVec_10_T_3[6:0] ? myVec_56 : _GEN_15201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15203 = 7'h39 == _myNewVec_10_T_3[6:0] ? myVec_57 : _GEN_15202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15204 = 7'h3a == _myNewVec_10_T_3[6:0] ? myVec_58 : _GEN_15203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15205 = 7'h3b == _myNewVec_10_T_3[6:0] ? myVec_59 : _GEN_15204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15206 = 7'h3c == _myNewVec_10_T_3[6:0] ? myVec_60 : _GEN_15205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15207 = 7'h3d == _myNewVec_10_T_3[6:0] ? myVec_61 : _GEN_15206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15208 = 7'h3e == _myNewVec_10_T_3[6:0] ? myVec_62 : _GEN_15207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15209 = 7'h3f == _myNewVec_10_T_3[6:0] ? myVec_63 : _GEN_15208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15210 = 7'h40 == _myNewVec_10_T_3[6:0] ? myVec_64 : _GEN_15209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15211 = 7'h41 == _myNewVec_10_T_3[6:0] ? myVec_65 : _GEN_15210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15212 = 7'h42 == _myNewVec_10_T_3[6:0] ? myVec_66 : _GEN_15211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15213 = 7'h43 == _myNewVec_10_T_3[6:0] ? myVec_67 : _GEN_15212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15214 = 7'h44 == _myNewVec_10_T_3[6:0] ? myVec_68 : _GEN_15213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15215 = 7'h45 == _myNewVec_10_T_3[6:0] ? myVec_69 : _GEN_15214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15216 = 7'h46 == _myNewVec_10_T_3[6:0] ? myVec_70 : _GEN_15215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15217 = 7'h47 == _myNewVec_10_T_3[6:0] ? myVec_71 : _GEN_15216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15218 = 7'h48 == _myNewVec_10_T_3[6:0] ? myVec_72 : _GEN_15217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15219 = 7'h49 == _myNewVec_10_T_3[6:0] ? myVec_73 : _GEN_15218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15220 = 7'h4a == _myNewVec_10_T_3[6:0] ? myVec_74 : _GEN_15219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15221 = 7'h4b == _myNewVec_10_T_3[6:0] ? myVec_75 : _GEN_15220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15222 = 7'h4c == _myNewVec_10_T_3[6:0] ? myVec_76 : _GEN_15221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15223 = 7'h4d == _myNewVec_10_T_3[6:0] ? myVec_77 : _GEN_15222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15224 = 7'h4e == _myNewVec_10_T_3[6:0] ? myVec_78 : _GEN_15223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15225 = 7'h4f == _myNewVec_10_T_3[6:0] ? myVec_79 : _GEN_15224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15226 = 7'h50 == _myNewVec_10_T_3[6:0] ? myVec_80 : _GEN_15225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15227 = 7'h51 == _myNewVec_10_T_3[6:0] ? myVec_81 : _GEN_15226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15228 = 7'h52 == _myNewVec_10_T_3[6:0] ? myVec_82 : _GEN_15227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15229 = 7'h53 == _myNewVec_10_T_3[6:0] ? myVec_83 : _GEN_15228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15230 = 7'h54 == _myNewVec_10_T_3[6:0] ? myVec_84 : _GEN_15229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15231 = 7'h55 == _myNewVec_10_T_3[6:0] ? myVec_85 : _GEN_15230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15232 = 7'h56 == _myNewVec_10_T_3[6:0] ? myVec_86 : _GEN_15231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15233 = 7'h57 == _myNewVec_10_T_3[6:0] ? myVec_87 : _GEN_15232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15234 = 7'h58 == _myNewVec_10_T_3[6:0] ? myVec_88 : _GEN_15233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15235 = 7'h59 == _myNewVec_10_T_3[6:0] ? myVec_89 : _GEN_15234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15236 = 7'h5a == _myNewVec_10_T_3[6:0] ? myVec_90 : _GEN_15235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15237 = 7'h5b == _myNewVec_10_T_3[6:0] ? myVec_91 : _GEN_15236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15238 = 7'h5c == _myNewVec_10_T_3[6:0] ? myVec_92 : _GEN_15237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15239 = 7'h5d == _myNewVec_10_T_3[6:0] ? myVec_93 : _GEN_15238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15240 = 7'h5e == _myNewVec_10_T_3[6:0] ? myVec_94 : _GEN_15239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15241 = 7'h5f == _myNewVec_10_T_3[6:0] ? myVec_95 : _GEN_15240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15242 = 7'h60 == _myNewVec_10_T_3[6:0] ? myVec_96 : _GEN_15241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15243 = 7'h61 == _myNewVec_10_T_3[6:0] ? myVec_97 : _GEN_15242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15244 = 7'h62 == _myNewVec_10_T_3[6:0] ? myVec_98 : _GEN_15243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15245 = 7'h63 == _myNewVec_10_T_3[6:0] ? myVec_99 : _GEN_15244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15246 = 7'h64 == _myNewVec_10_T_3[6:0] ? myVec_100 : _GEN_15245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15247 = 7'h65 == _myNewVec_10_T_3[6:0] ? myVec_101 : _GEN_15246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15248 = 7'h66 == _myNewVec_10_T_3[6:0] ? myVec_102 : _GEN_15247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15249 = 7'h67 == _myNewVec_10_T_3[6:0] ? myVec_103 : _GEN_15248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15250 = 7'h68 == _myNewVec_10_T_3[6:0] ? myVec_104 : _GEN_15249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15251 = 7'h69 == _myNewVec_10_T_3[6:0] ? myVec_105 : _GEN_15250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15252 = 7'h6a == _myNewVec_10_T_3[6:0] ? myVec_106 : _GEN_15251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15253 = 7'h6b == _myNewVec_10_T_3[6:0] ? myVec_107 : _GEN_15252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15254 = 7'h6c == _myNewVec_10_T_3[6:0] ? myVec_108 : _GEN_15253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15255 = 7'h6d == _myNewVec_10_T_3[6:0] ? myVec_109 : _GEN_15254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15256 = 7'h6e == _myNewVec_10_T_3[6:0] ? myVec_110 : _GEN_15255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15257 = 7'h6f == _myNewVec_10_T_3[6:0] ? myVec_111 : _GEN_15256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15258 = 7'h70 == _myNewVec_10_T_3[6:0] ? myVec_112 : _GEN_15257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15259 = 7'h71 == _myNewVec_10_T_3[6:0] ? myVec_113 : _GEN_15258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15260 = 7'h72 == _myNewVec_10_T_3[6:0] ? myVec_114 : _GEN_15259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15261 = 7'h73 == _myNewVec_10_T_3[6:0] ? myVec_115 : _GEN_15260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15262 = 7'h74 == _myNewVec_10_T_3[6:0] ? myVec_116 : _GEN_15261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15263 = 7'h75 == _myNewVec_10_T_3[6:0] ? myVec_117 : _GEN_15262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15264 = 7'h76 == _myNewVec_10_T_3[6:0] ? myVec_118 : _GEN_15263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15265 = 7'h77 == _myNewVec_10_T_3[6:0] ? myVec_119 : _GEN_15264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15266 = 7'h78 == _myNewVec_10_T_3[6:0] ? myVec_120 : _GEN_15265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15267 = 7'h79 == _myNewVec_10_T_3[6:0] ? myVec_121 : _GEN_15266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15268 = 7'h7a == _myNewVec_10_T_3[6:0] ? myVec_122 : _GEN_15267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15269 = 7'h7b == _myNewVec_10_T_3[6:0] ? myVec_123 : _GEN_15268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15270 = 7'h7c == _myNewVec_10_T_3[6:0] ? myVec_124 : _GEN_15269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15271 = 7'h7d == _myNewVec_10_T_3[6:0] ? myVec_125 : _GEN_15270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15272 = 7'h7e == _myNewVec_10_T_3[6:0] ? myVec_126 : _GEN_15271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_10 = 7'h7f == _myNewVec_10_T_3[6:0] ? myVec_127 : _GEN_15272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_9_T_3 = _myNewVec_127_T_1 + 16'h76; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_15275 = 7'h1 == _myNewVec_9_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15276 = 7'h2 == _myNewVec_9_T_3[6:0] ? myVec_2 : _GEN_15275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15277 = 7'h3 == _myNewVec_9_T_3[6:0] ? myVec_3 : _GEN_15276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15278 = 7'h4 == _myNewVec_9_T_3[6:0] ? myVec_4 : _GEN_15277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15279 = 7'h5 == _myNewVec_9_T_3[6:0] ? myVec_5 : _GEN_15278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15280 = 7'h6 == _myNewVec_9_T_3[6:0] ? myVec_6 : _GEN_15279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15281 = 7'h7 == _myNewVec_9_T_3[6:0] ? myVec_7 : _GEN_15280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15282 = 7'h8 == _myNewVec_9_T_3[6:0] ? myVec_8 : _GEN_15281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15283 = 7'h9 == _myNewVec_9_T_3[6:0] ? myVec_9 : _GEN_15282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15284 = 7'ha == _myNewVec_9_T_3[6:0] ? myVec_10 : _GEN_15283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15285 = 7'hb == _myNewVec_9_T_3[6:0] ? myVec_11 : _GEN_15284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15286 = 7'hc == _myNewVec_9_T_3[6:0] ? myVec_12 : _GEN_15285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15287 = 7'hd == _myNewVec_9_T_3[6:0] ? myVec_13 : _GEN_15286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15288 = 7'he == _myNewVec_9_T_3[6:0] ? myVec_14 : _GEN_15287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15289 = 7'hf == _myNewVec_9_T_3[6:0] ? myVec_15 : _GEN_15288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15290 = 7'h10 == _myNewVec_9_T_3[6:0] ? myVec_16 : _GEN_15289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15291 = 7'h11 == _myNewVec_9_T_3[6:0] ? myVec_17 : _GEN_15290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15292 = 7'h12 == _myNewVec_9_T_3[6:0] ? myVec_18 : _GEN_15291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15293 = 7'h13 == _myNewVec_9_T_3[6:0] ? myVec_19 : _GEN_15292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15294 = 7'h14 == _myNewVec_9_T_3[6:0] ? myVec_20 : _GEN_15293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15295 = 7'h15 == _myNewVec_9_T_3[6:0] ? myVec_21 : _GEN_15294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15296 = 7'h16 == _myNewVec_9_T_3[6:0] ? myVec_22 : _GEN_15295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15297 = 7'h17 == _myNewVec_9_T_3[6:0] ? myVec_23 : _GEN_15296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15298 = 7'h18 == _myNewVec_9_T_3[6:0] ? myVec_24 : _GEN_15297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15299 = 7'h19 == _myNewVec_9_T_3[6:0] ? myVec_25 : _GEN_15298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15300 = 7'h1a == _myNewVec_9_T_3[6:0] ? myVec_26 : _GEN_15299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15301 = 7'h1b == _myNewVec_9_T_3[6:0] ? myVec_27 : _GEN_15300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15302 = 7'h1c == _myNewVec_9_T_3[6:0] ? myVec_28 : _GEN_15301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15303 = 7'h1d == _myNewVec_9_T_3[6:0] ? myVec_29 : _GEN_15302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15304 = 7'h1e == _myNewVec_9_T_3[6:0] ? myVec_30 : _GEN_15303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15305 = 7'h1f == _myNewVec_9_T_3[6:0] ? myVec_31 : _GEN_15304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15306 = 7'h20 == _myNewVec_9_T_3[6:0] ? myVec_32 : _GEN_15305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15307 = 7'h21 == _myNewVec_9_T_3[6:0] ? myVec_33 : _GEN_15306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15308 = 7'h22 == _myNewVec_9_T_3[6:0] ? myVec_34 : _GEN_15307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15309 = 7'h23 == _myNewVec_9_T_3[6:0] ? myVec_35 : _GEN_15308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15310 = 7'h24 == _myNewVec_9_T_3[6:0] ? myVec_36 : _GEN_15309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15311 = 7'h25 == _myNewVec_9_T_3[6:0] ? myVec_37 : _GEN_15310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15312 = 7'h26 == _myNewVec_9_T_3[6:0] ? myVec_38 : _GEN_15311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15313 = 7'h27 == _myNewVec_9_T_3[6:0] ? myVec_39 : _GEN_15312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15314 = 7'h28 == _myNewVec_9_T_3[6:0] ? myVec_40 : _GEN_15313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15315 = 7'h29 == _myNewVec_9_T_3[6:0] ? myVec_41 : _GEN_15314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15316 = 7'h2a == _myNewVec_9_T_3[6:0] ? myVec_42 : _GEN_15315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15317 = 7'h2b == _myNewVec_9_T_3[6:0] ? myVec_43 : _GEN_15316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15318 = 7'h2c == _myNewVec_9_T_3[6:0] ? myVec_44 : _GEN_15317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15319 = 7'h2d == _myNewVec_9_T_3[6:0] ? myVec_45 : _GEN_15318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15320 = 7'h2e == _myNewVec_9_T_3[6:0] ? myVec_46 : _GEN_15319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15321 = 7'h2f == _myNewVec_9_T_3[6:0] ? myVec_47 : _GEN_15320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15322 = 7'h30 == _myNewVec_9_T_3[6:0] ? myVec_48 : _GEN_15321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15323 = 7'h31 == _myNewVec_9_T_3[6:0] ? myVec_49 : _GEN_15322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15324 = 7'h32 == _myNewVec_9_T_3[6:0] ? myVec_50 : _GEN_15323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15325 = 7'h33 == _myNewVec_9_T_3[6:0] ? myVec_51 : _GEN_15324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15326 = 7'h34 == _myNewVec_9_T_3[6:0] ? myVec_52 : _GEN_15325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15327 = 7'h35 == _myNewVec_9_T_3[6:0] ? myVec_53 : _GEN_15326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15328 = 7'h36 == _myNewVec_9_T_3[6:0] ? myVec_54 : _GEN_15327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15329 = 7'h37 == _myNewVec_9_T_3[6:0] ? myVec_55 : _GEN_15328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15330 = 7'h38 == _myNewVec_9_T_3[6:0] ? myVec_56 : _GEN_15329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15331 = 7'h39 == _myNewVec_9_T_3[6:0] ? myVec_57 : _GEN_15330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15332 = 7'h3a == _myNewVec_9_T_3[6:0] ? myVec_58 : _GEN_15331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15333 = 7'h3b == _myNewVec_9_T_3[6:0] ? myVec_59 : _GEN_15332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15334 = 7'h3c == _myNewVec_9_T_3[6:0] ? myVec_60 : _GEN_15333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15335 = 7'h3d == _myNewVec_9_T_3[6:0] ? myVec_61 : _GEN_15334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15336 = 7'h3e == _myNewVec_9_T_3[6:0] ? myVec_62 : _GEN_15335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15337 = 7'h3f == _myNewVec_9_T_3[6:0] ? myVec_63 : _GEN_15336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15338 = 7'h40 == _myNewVec_9_T_3[6:0] ? myVec_64 : _GEN_15337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15339 = 7'h41 == _myNewVec_9_T_3[6:0] ? myVec_65 : _GEN_15338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15340 = 7'h42 == _myNewVec_9_T_3[6:0] ? myVec_66 : _GEN_15339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15341 = 7'h43 == _myNewVec_9_T_3[6:0] ? myVec_67 : _GEN_15340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15342 = 7'h44 == _myNewVec_9_T_3[6:0] ? myVec_68 : _GEN_15341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15343 = 7'h45 == _myNewVec_9_T_3[6:0] ? myVec_69 : _GEN_15342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15344 = 7'h46 == _myNewVec_9_T_3[6:0] ? myVec_70 : _GEN_15343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15345 = 7'h47 == _myNewVec_9_T_3[6:0] ? myVec_71 : _GEN_15344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15346 = 7'h48 == _myNewVec_9_T_3[6:0] ? myVec_72 : _GEN_15345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15347 = 7'h49 == _myNewVec_9_T_3[6:0] ? myVec_73 : _GEN_15346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15348 = 7'h4a == _myNewVec_9_T_3[6:0] ? myVec_74 : _GEN_15347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15349 = 7'h4b == _myNewVec_9_T_3[6:0] ? myVec_75 : _GEN_15348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15350 = 7'h4c == _myNewVec_9_T_3[6:0] ? myVec_76 : _GEN_15349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15351 = 7'h4d == _myNewVec_9_T_3[6:0] ? myVec_77 : _GEN_15350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15352 = 7'h4e == _myNewVec_9_T_3[6:0] ? myVec_78 : _GEN_15351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15353 = 7'h4f == _myNewVec_9_T_3[6:0] ? myVec_79 : _GEN_15352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15354 = 7'h50 == _myNewVec_9_T_3[6:0] ? myVec_80 : _GEN_15353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15355 = 7'h51 == _myNewVec_9_T_3[6:0] ? myVec_81 : _GEN_15354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15356 = 7'h52 == _myNewVec_9_T_3[6:0] ? myVec_82 : _GEN_15355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15357 = 7'h53 == _myNewVec_9_T_3[6:0] ? myVec_83 : _GEN_15356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15358 = 7'h54 == _myNewVec_9_T_3[6:0] ? myVec_84 : _GEN_15357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15359 = 7'h55 == _myNewVec_9_T_3[6:0] ? myVec_85 : _GEN_15358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15360 = 7'h56 == _myNewVec_9_T_3[6:0] ? myVec_86 : _GEN_15359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15361 = 7'h57 == _myNewVec_9_T_3[6:0] ? myVec_87 : _GEN_15360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15362 = 7'h58 == _myNewVec_9_T_3[6:0] ? myVec_88 : _GEN_15361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15363 = 7'h59 == _myNewVec_9_T_3[6:0] ? myVec_89 : _GEN_15362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15364 = 7'h5a == _myNewVec_9_T_3[6:0] ? myVec_90 : _GEN_15363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15365 = 7'h5b == _myNewVec_9_T_3[6:0] ? myVec_91 : _GEN_15364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15366 = 7'h5c == _myNewVec_9_T_3[6:0] ? myVec_92 : _GEN_15365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15367 = 7'h5d == _myNewVec_9_T_3[6:0] ? myVec_93 : _GEN_15366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15368 = 7'h5e == _myNewVec_9_T_3[6:0] ? myVec_94 : _GEN_15367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15369 = 7'h5f == _myNewVec_9_T_3[6:0] ? myVec_95 : _GEN_15368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15370 = 7'h60 == _myNewVec_9_T_3[6:0] ? myVec_96 : _GEN_15369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15371 = 7'h61 == _myNewVec_9_T_3[6:0] ? myVec_97 : _GEN_15370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15372 = 7'h62 == _myNewVec_9_T_3[6:0] ? myVec_98 : _GEN_15371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15373 = 7'h63 == _myNewVec_9_T_3[6:0] ? myVec_99 : _GEN_15372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15374 = 7'h64 == _myNewVec_9_T_3[6:0] ? myVec_100 : _GEN_15373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15375 = 7'h65 == _myNewVec_9_T_3[6:0] ? myVec_101 : _GEN_15374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15376 = 7'h66 == _myNewVec_9_T_3[6:0] ? myVec_102 : _GEN_15375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15377 = 7'h67 == _myNewVec_9_T_3[6:0] ? myVec_103 : _GEN_15376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15378 = 7'h68 == _myNewVec_9_T_3[6:0] ? myVec_104 : _GEN_15377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15379 = 7'h69 == _myNewVec_9_T_3[6:0] ? myVec_105 : _GEN_15378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15380 = 7'h6a == _myNewVec_9_T_3[6:0] ? myVec_106 : _GEN_15379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15381 = 7'h6b == _myNewVec_9_T_3[6:0] ? myVec_107 : _GEN_15380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15382 = 7'h6c == _myNewVec_9_T_3[6:0] ? myVec_108 : _GEN_15381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15383 = 7'h6d == _myNewVec_9_T_3[6:0] ? myVec_109 : _GEN_15382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15384 = 7'h6e == _myNewVec_9_T_3[6:0] ? myVec_110 : _GEN_15383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15385 = 7'h6f == _myNewVec_9_T_3[6:0] ? myVec_111 : _GEN_15384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15386 = 7'h70 == _myNewVec_9_T_3[6:0] ? myVec_112 : _GEN_15385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15387 = 7'h71 == _myNewVec_9_T_3[6:0] ? myVec_113 : _GEN_15386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15388 = 7'h72 == _myNewVec_9_T_3[6:0] ? myVec_114 : _GEN_15387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15389 = 7'h73 == _myNewVec_9_T_3[6:0] ? myVec_115 : _GEN_15388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15390 = 7'h74 == _myNewVec_9_T_3[6:0] ? myVec_116 : _GEN_15389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15391 = 7'h75 == _myNewVec_9_T_3[6:0] ? myVec_117 : _GEN_15390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15392 = 7'h76 == _myNewVec_9_T_3[6:0] ? myVec_118 : _GEN_15391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15393 = 7'h77 == _myNewVec_9_T_3[6:0] ? myVec_119 : _GEN_15392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15394 = 7'h78 == _myNewVec_9_T_3[6:0] ? myVec_120 : _GEN_15393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15395 = 7'h79 == _myNewVec_9_T_3[6:0] ? myVec_121 : _GEN_15394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15396 = 7'h7a == _myNewVec_9_T_3[6:0] ? myVec_122 : _GEN_15395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15397 = 7'h7b == _myNewVec_9_T_3[6:0] ? myVec_123 : _GEN_15396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15398 = 7'h7c == _myNewVec_9_T_3[6:0] ? myVec_124 : _GEN_15397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15399 = 7'h7d == _myNewVec_9_T_3[6:0] ? myVec_125 : _GEN_15398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15400 = 7'h7e == _myNewVec_9_T_3[6:0] ? myVec_126 : _GEN_15399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_9 = 7'h7f == _myNewVec_9_T_3[6:0] ? myVec_127 : _GEN_15400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_8_T_3 = _myNewVec_127_T_1 + 16'h77; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_15403 = 7'h1 == _myNewVec_8_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15404 = 7'h2 == _myNewVec_8_T_3[6:0] ? myVec_2 : _GEN_15403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15405 = 7'h3 == _myNewVec_8_T_3[6:0] ? myVec_3 : _GEN_15404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15406 = 7'h4 == _myNewVec_8_T_3[6:0] ? myVec_4 : _GEN_15405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15407 = 7'h5 == _myNewVec_8_T_3[6:0] ? myVec_5 : _GEN_15406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15408 = 7'h6 == _myNewVec_8_T_3[6:0] ? myVec_6 : _GEN_15407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15409 = 7'h7 == _myNewVec_8_T_3[6:0] ? myVec_7 : _GEN_15408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15410 = 7'h8 == _myNewVec_8_T_3[6:0] ? myVec_8 : _GEN_15409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15411 = 7'h9 == _myNewVec_8_T_3[6:0] ? myVec_9 : _GEN_15410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15412 = 7'ha == _myNewVec_8_T_3[6:0] ? myVec_10 : _GEN_15411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15413 = 7'hb == _myNewVec_8_T_3[6:0] ? myVec_11 : _GEN_15412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15414 = 7'hc == _myNewVec_8_T_3[6:0] ? myVec_12 : _GEN_15413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15415 = 7'hd == _myNewVec_8_T_3[6:0] ? myVec_13 : _GEN_15414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15416 = 7'he == _myNewVec_8_T_3[6:0] ? myVec_14 : _GEN_15415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15417 = 7'hf == _myNewVec_8_T_3[6:0] ? myVec_15 : _GEN_15416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15418 = 7'h10 == _myNewVec_8_T_3[6:0] ? myVec_16 : _GEN_15417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15419 = 7'h11 == _myNewVec_8_T_3[6:0] ? myVec_17 : _GEN_15418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15420 = 7'h12 == _myNewVec_8_T_3[6:0] ? myVec_18 : _GEN_15419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15421 = 7'h13 == _myNewVec_8_T_3[6:0] ? myVec_19 : _GEN_15420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15422 = 7'h14 == _myNewVec_8_T_3[6:0] ? myVec_20 : _GEN_15421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15423 = 7'h15 == _myNewVec_8_T_3[6:0] ? myVec_21 : _GEN_15422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15424 = 7'h16 == _myNewVec_8_T_3[6:0] ? myVec_22 : _GEN_15423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15425 = 7'h17 == _myNewVec_8_T_3[6:0] ? myVec_23 : _GEN_15424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15426 = 7'h18 == _myNewVec_8_T_3[6:0] ? myVec_24 : _GEN_15425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15427 = 7'h19 == _myNewVec_8_T_3[6:0] ? myVec_25 : _GEN_15426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15428 = 7'h1a == _myNewVec_8_T_3[6:0] ? myVec_26 : _GEN_15427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15429 = 7'h1b == _myNewVec_8_T_3[6:0] ? myVec_27 : _GEN_15428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15430 = 7'h1c == _myNewVec_8_T_3[6:0] ? myVec_28 : _GEN_15429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15431 = 7'h1d == _myNewVec_8_T_3[6:0] ? myVec_29 : _GEN_15430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15432 = 7'h1e == _myNewVec_8_T_3[6:0] ? myVec_30 : _GEN_15431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15433 = 7'h1f == _myNewVec_8_T_3[6:0] ? myVec_31 : _GEN_15432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15434 = 7'h20 == _myNewVec_8_T_3[6:0] ? myVec_32 : _GEN_15433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15435 = 7'h21 == _myNewVec_8_T_3[6:0] ? myVec_33 : _GEN_15434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15436 = 7'h22 == _myNewVec_8_T_3[6:0] ? myVec_34 : _GEN_15435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15437 = 7'h23 == _myNewVec_8_T_3[6:0] ? myVec_35 : _GEN_15436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15438 = 7'h24 == _myNewVec_8_T_3[6:0] ? myVec_36 : _GEN_15437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15439 = 7'h25 == _myNewVec_8_T_3[6:0] ? myVec_37 : _GEN_15438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15440 = 7'h26 == _myNewVec_8_T_3[6:0] ? myVec_38 : _GEN_15439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15441 = 7'h27 == _myNewVec_8_T_3[6:0] ? myVec_39 : _GEN_15440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15442 = 7'h28 == _myNewVec_8_T_3[6:0] ? myVec_40 : _GEN_15441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15443 = 7'h29 == _myNewVec_8_T_3[6:0] ? myVec_41 : _GEN_15442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15444 = 7'h2a == _myNewVec_8_T_3[6:0] ? myVec_42 : _GEN_15443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15445 = 7'h2b == _myNewVec_8_T_3[6:0] ? myVec_43 : _GEN_15444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15446 = 7'h2c == _myNewVec_8_T_3[6:0] ? myVec_44 : _GEN_15445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15447 = 7'h2d == _myNewVec_8_T_3[6:0] ? myVec_45 : _GEN_15446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15448 = 7'h2e == _myNewVec_8_T_3[6:0] ? myVec_46 : _GEN_15447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15449 = 7'h2f == _myNewVec_8_T_3[6:0] ? myVec_47 : _GEN_15448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15450 = 7'h30 == _myNewVec_8_T_3[6:0] ? myVec_48 : _GEN_15449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15451 = 7'h31 == _myNewVec_8_T_3[6:0] ? myVec_49 : _GEN_15450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15452 = 7'h32 == _myNewVec_8_T_3[6:0] ? myVec_50 : _GEN_15451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15453 = 7'h33 == _myNewVec_8_T_3[6:0] ? myVec_51 : _GEN_15452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15454 = 7'h34 == _myNewVec_8_T_3[6:0] ? myVec_52 : _GEN_15453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15455 = 7'h35 == _myNewVec_8_T_3[6:0] ? myVec_53 : _GEN_15454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15456 = 7'h36 == _myNewVec_8_T_3[6:0] ? myVec_54 : _GEN_15455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15457 = 7'h37 == _myNewVec_8_T_3[6:0] ? myVec_55 : _GEN_15456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15458 = 7'h38 == _myNewVec_8_T_3[6:0] ? myVec_56 : _GEN_15457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15459 = 7'h39 == _myNewVec_8_T_3[6:0] ? myVec_57 : _GEN_15458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15460 = 7'h3a == _myNewVec_8_T_3[6:0] ? myVec_58 : _GEN_15459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15461 = 7'h3b == _myNewVec_8_T_3[6:0] ? myVec_59 : _GEN_15460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15462 = 7'h3c == _myNewVec_8_T_3[6:0] ? myVec_60 : _GEN_15461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15463 = 7'h3d == _myNewVec_8_T_3[6:0] ? myVec_61 : _GEN_15462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15464 = 7'h3e == _myNewVec_8_T_3[6:0] ? myVec_62 : _GEN_15463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15465 = 7'h3f == _myNewVec_8_T_3[6:0] ? myVec_63 : _GEN_15464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15466 = 7'h40 == _myNewVec_8_T_3[6:0] ? myVec_64 : _GEN_15465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15467 = 7'h41 == _myNewVec_8_T_3[6:0] ? myVec_65 : _GEN_15466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15468 = 7'h42 == _myNewVec_8_T_3[6:0] ? myVec_66 : _GEN_15467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15469 = 7'h43 == _myNewVec_8_T_3[6:0] ? myVec_67 : _GEN_15468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15470 = 7'h44 == _myNewVec_8_T_3[6:0] ? myVec_68 : _GEN_15469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15471 = 7'h45 == _myNewVec_8_T_3[6:0] ? myVec_69 : _GEN_15470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15472 = 7'h46 == _myNewVec_8_T_3[6:0] ? myVec_70 : _GEN_15471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15473 = 7'h47 == _myNewVec_8_T_3[6:0] ? myVec_71 : _GEN_15472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15474 = 7'h48 == _myNewVec_8_T_3[6:0] ? myVec_72 : _GEN_15473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15475 = 7'h49 == _myNewVec_8_T_3[6:0] ? myVec_73 : _GEN_15474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15476 = 7'h4a == _myNewVec_8_T_3[6:0] ? myVec_74 : _GEN_15475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15477 = 7'h4b == _myNewVec_8_T_3[6:0] ? myVec_75 : _GEN_15476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15478 = 7'h4c == _myNewVec_8_T_3[6:0] ? myVec_76 : _GEN_15477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15479 = 7'h4d == _myNewVec_8_T_3[6:0] ? myVec_77 : _GEN_15478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15480 = 7'h4e == _myNewVec_8_T_3[6:0] ? myVec_78 : _GEN_15479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15481 = 7'h4f == _myNewVec_8_T_3[6:0] ? myVec_79 : _GEN_15480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15482 = 7'h50 == _myNewVec_8_T_3[6:0] ? myVec_80 : _GEN_15481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15483 = 7'h51 == _myNewVec_8_T_3[6:0] ? myVec_81 : _GEN_15482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15484 = 7'h52 == _myNewVec_8_T_3[6:0] ? myVec_82 : _GEN_15483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15485 = 7'h53 == _myNewVec_8_T_3[6:0] ? myVec_83 : _GEN_15484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15486 = 7'h54 == _myNewVec_8_T_3[6:0] ? myVec_84 : _GEN_15485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15487 = 7'h55 == _myNewVec_8_T_3[6:0] ? myVec_85 : _GEN_15486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15488 = 7'h56 == _myNewVec_8_T_3[6:0] ? myVec_86 : _GEN_15487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15489 = 7'h57 == _myNewVec_8_T_3[6:0] ? myVec_87 : _GEN_15488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15490 = 7'h58 == _myNewVec_8_T_3[6:0] ? myVec_88 : _GEN_15489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15491 = 7'h59 == _myNewVec_8_T_3[6:0] ? myVec_89 : _GEN_15490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15492 = 7'h5a == _myNewVec_8_T_3[6:0] ? myVec_90 : _GEN_15491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15493 = 7'h5b == _myNewVec_8_T_3[6:0] ? myVec_91 : _GEN_15492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15494 = 7'h5c == _myNewVec_8_T_3[6:0] ? myVec_92 : _GEN_15493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15495 = 7'h5d == _myNewVec_8_T_3[6:0] ? myVec_93 : _GEN_15494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15496 = 7'h5e == _myNewVec_8_T_3[6:0] ? myVec_94 : _GEN_15495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15497 = 7'h5f == _myNewVec_8_T_3[6:0] ? myVec_95 : _GEN_15496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15498 = 7'h60 == _myNewVec_8_T_3[6:0] ? myVec_96 : _GEN_15497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15499 = 7'h61 == _myNewVec_8_T_3[6:0] ? myVec_97 : _GEN_15498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15500 = 7'h62 == _myNewVec_8_T_3[6:0] ? myVec_98 : _GEN_15499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15501 = 7'h63 == _myNewVec_8_T_3[6:0] ? myVec_99 : _GEN_15500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15502 = 7'h64 == _myNewVec_8_T_3[6:0] ? myVec_100 : _GEN_15501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15503 = 7'h65 == _myNewVec_8_T_3[6:0] ? myVec_101 : _GEN_15502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15504 = 7'h66 == _myNewVec_8_T_3[6:0] ? myVec_102 : _GEN_15503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15505 = 7'h67 == _myNewVec_8_T_3[6:0] ? myVec_103 : _GEN_15504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15506 = 7'h68 == _myNewVec_8_T_3[6:0] ? myVec_104 : _GEN_15505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15507 = 7'h69 == _myNewVec_8_T_3[6:0] ? myVec_105 : _GEN_15506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15508 = 7'h6a == _myNewVec_8_T_3[6:0] ? myVec_106 : _GEN_15507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15509 = 7'h6b == _myNewVec_8_T_3[6:0] ? myVec_107 : _GEN_15508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15510 = 7'h6c == _myNewVec_8_T_3[6:0] ? myVec_108 : _GEN_15509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15511 = 7'h6d == _myNewVec_8_T_3[6:0] ? myVec_109 : _GEN_15510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15512 = 7'h6e == _myNewVec_8_T_3[6:0] ? myVec_110 : _GEN_15511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15513 = 7'h6f == _myNewVec_8_T_3[6:0] ? myVec_111 : _GEN_15512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15514 = 7'h70 == _myNewVec_8_T_3[6:0] ? myVec_112 : _GEN_15513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15515 = 7'h71 == _myNewVec_8_T_3[6:0] ? myVec_113 : _GEN_15514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15516 = 7'h72 == _myNewVec_8_T_3[6:0] ? myVec_114 : _GEN_15515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15517 = 7'h73 == _myNewVec_8_T_3[6:0] ? myVec_115 : _GEN_15516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15518 = 7'h74 == _myNewVec_8_T_3[6:0] ? myVec_116 : _GEN_15517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15519 = 7'h75 == _myNewVec_8_T_3[6:0] ? myVec_117 : _GEN_15518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15520 = 7'h76 == _myNewVec_8_T_3[6:0] ? myVec_118 : _GEN_15519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15521 = 7'h77 == _myNewVec_8_T_3[6:0] ? myVec_119 : _GEN_15520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15522 = 7'h78 == _myNewVec_8_T_3[6:0] ? myVec_120 : _GEN_15521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15523 = 7'h79 == _myNewVec_8_T_3[6:0] ? myVec_121 : _GEN_15522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15524 = 7'h7a == _myNewVec_8_T_3[6:0] ? myVec_122 : _GEN_15523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15525 = 7'h7b == _myNewVec_8_T_3[6:0] ? myVec_123 : _GEN_15524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15526 = 7'h7c == _myNewVec_8_T_3[6:0] ? myVec_124 : _GEN_15525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15527 = 7'h7d == _myNewVec_8_T_3[6:0] ? myVec_125 : _GEN_15526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15528 = 7'h7e == _myNewVec_8_T_3[6:0] ? myVec_126 : _GEN_15527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_8 = 7'h7f == _myNewVec_8_T_3[6:0] ? myVec_127 : _GEN_15528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_7_T_3 = _myNewVec_127_T_1 + 16'h78; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_15531 = 7'h1 == _myNewVec_7_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15532 = 7'h2 == _myNewVec_7_T_3[6:0] ? myVec_2 : _GEN_15531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15533 = 7'h3 == _myNewVec_7_T_3[6:0] ? myVec_3 : _GEN_15532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15534 = 7'h4 == _myNewVec_7_T_3[6:0] ? myVec_4 : _GEN_15533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15535 = 7'h5 == _myNewVec_7_T_3[6:0] ? myVec_5 : _GEN_15534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15536 = 7'h6 == _myNewVec_7_T_3[6:0] ? myVec_6 : _GEN_15535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15537 = 7'h7 == _myNewVec_7_T_3[6:0] ? myVec_7 : _GEN_15536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15538 = 7'h8 == _myNewVec_7_T_3[6:0] ? myVec_8 : _GEN_15537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15539 = 7'h9 == _myNewVec_7_T_3[6:0] ? myVec_9 : _GEN_15538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15540 = 7'ha == _myNewVec_7_T_3[6:0] ? myVec_10 : _GEN_15539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15541 = 7'hb == _myNewVec_7_T_3[6:0] ? myVec_11 : _GEN_15540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15542 = 7'hc == _myNewVec_7_T_3[6:0] ? myVec_12 : _GEN_15541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15543 = 7'hd == _myNewVec_7_T_3[6:0] ? myVec_13 : _GEN_15542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15544 = 7'he == _myNewVec_7_T_3[6:0] ? myVec_14 : _GEN_15543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15545 = 7'hf == _myNewVec_7_T_3[6:0] ? myVec_15 : _GEN_15544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15546 = 7'h10 == _myNewVec_7_T_3[6:0] ? myVec_16 : _GEN_15545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15547 = 7'h11 == _myNewVec_7_T_3[6:0] ? myVec_17 : _GEN_15546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15548 = 7'h12 == _myNewVec_7_T_3[6:0] ? myVec_18 : _GEN_15547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15549 = 7'h13 == _myNewVec_7_T_3[6:0] ? myVec_19 : _GEN_15548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15550 = 7'h14 == _myNewVec_7_T_3[6:0] ? myVec_20 : _GEN_15549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15551 = 7'h15 == _myNewVec_7_T_3[6:0] ? myVec_21 : _GEN_15550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15552 = 7'h16 == _myNewVec_7_T_3[6:0] ? myVec_22 : _GEN_15551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15553 = 7'h17 == _myNewVec_7_T_3[6:0] ? myVec_23 : _GEN_15552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15554 = 7'h18 == _myNewVec_7_T_3[6:0] ? myVec_24 : _GEN_15553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15555 = 7'h19 == _myNewVec_7_T_3[6:0] ? myVec_25 : _GEN_15554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15556 = 7'h1a == _myNewVec_7_T_3[6:0] ? myVec_26 : _GEN_15555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15557 = 7'h1b == _myNewVec_7_T_3[6:0] ? myVec_27 : _GEN_15556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15558 = 7'h1c == _myNewVec_7_T_3[6:0] ? myVec_28 : _GEN_15557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15559 = 7'h1d == _myNewVec_7_T_3[6:0] ? myVec_29 : _GEN_15558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15560 = 7'h1e == _myNewVec_7_T_3[6:0] ? myVec_30 : _GEN_15559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15561 = 7'h1f == _myNewVec_7_T_3[6:0] ? myVec_31 : _GEN_15560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15562 = 7'h20 == _myNewVec_7_T_3[6:0] ? myVec_32 : _GEN_15561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15563 = 7'h21 == _myNewVec_7_T_3[6:0] ? myVec_33 : _GEN_15562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15564 = 7'h22 == _myNewVec_7_T_3[6:0] ? myVec_34 : _GEN_15563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15565 = 7'h23 == _myNewVec_7_T_3[6:0] ? myVec_35 : _GEN_15564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15566 = 7'h24 == _myNewVec_7_T_3[6:0] ? myVec_36 : _GEN_15565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15567 = 7'h25 == _myNewVec_7_T_3[6:0] ? myVec_37 : _GEN_15566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15568 = 7'h26 == _myNewVec_7_T_3[6:0] ? myVec_38 : _GEN_15567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15569 = 7'h27 == _myNewVec_7_T_3[6:0] ? myVec_39 : _GEN_15568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15570 = 7'h28 == _myNewVec_7_T_3[6:0] ? myVec_40 : _GEN_15569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15571 = 7'h29 == _myNewVec_7_T_3[6:0] ? myVec_41 : _GEN_15570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15572 = 7'h2a == _myNewVec_7_T_3[6:0] ? myVec_42 : _GEN_15571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15573 = 7'h2b == _myNewVec_7_T_3[6:0] ? myVec_43 : _GEN_15572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15574 = 7'h2c == _myNewVec_7_T_3[6:0] ? myVec_44 : _GEN_15573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15575 = 7'h2d == _myNewVec_7_T_3[6:0] ? myVec_45 : _GEN_15574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15576 = 7'h2e == _myNewVec_7_T_3[6:0] ? myVec_46 : _GEN_15575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15577 = 7'h2f == _myNewVec_7_T_3[6:0] ? myVec_47 : _GEN_15576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15578 = 7'h30 == _myNewVec_7_T_3[6:0] ? myVec_48 : _GEN_15577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15579 = 7'h31 == _myNewVec_7_T_3[6:0] ? myVec_49 : _GEN_15578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15580 = 7'h32 == _myNewVec_7_T_3[6:0] ? myVec_50 : _GEN_15579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15581 = 7'h33 == _myNewVec_7_T_3[6:0] ? myVec_51 : _GEN_15580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15582 = 7'h34 == _myNewVec_7_T_3[6:0] ? myVec_52 : _GEN_15581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15583 = 7'h35 == _myNewVec_7_T_3[6:0] ? myVec_53 : _GEN_15582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15584 = 7'h36 == _myNewVec_7_T_3[6:0] ? myVec_54 : _GEN_15583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15585 = 7'h37 == _myNewVec_7_T_3[6:0] ? myVec_55 : _GEN_15584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15586 = 7'h38 == _myNewVec_7_T_3[6:0] ? myVec_56 : _GEN_15585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15587 = 7'h39 == _myNewVec_7_T_3[6:0] ? myVec_57 : _GEN_15586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15588 = 7'h3a == _myNewVec_7_T_3[6:0] ? myVec_58 : _GEN_15587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15589 = 7'h3b == _myNewVec_7_T_3[6:0] ? myVec_59 : _GEN_15588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15590 = 7'h3c == _myNewVec_7_T_3[6:0] ? myVec_60 : _GEN_15589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15591 = 7'h3d == _myNewVec_7_T_3[6:0] ? myVec_61 : _GEN_15590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15592 = 7'h3e == _myNewVec_7_T_3[6:0] ? myVec_62 : _GEN_15591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15593 = 7'h3f == _myNewVec_7_T_3[6:0] ? myVec_63 : _GEN_15592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15594 = 7'h40 == _myNewVec_7_T_3[6:0] ? myVec_64 : _GEN_15593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15595 = 7'h41 == _myNewVec_7_T_3[6:0] ? myVec_65 : _GEN_15594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15596 = 7'h42 == _myNewVec_7_T_3[6:0] ? myVec_66 : _GEN_15595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15597 = 7'h43 == _myNewVec_7_T_3[6:0] ? myVec_67 : _GEN_15596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15598 = 7'h44 == _myNewVec_7_T_3[6:0] ? myVec_68 : _GEN_15597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15599 = 7'h45 == _myNewVec_7_T_3[6:0] ? myVec_69 : _GEN_15598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15600 = 7'h46 == _myNewVec_7_T_3[6:0] ? myVec_70 : _GEN_15599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15601 = 7'h47 == _myNewVec_7_T_3[6:0] ? myVec_71 : _GEN_15600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15602 = 7'h48 == _myNewVec_7_T_3[6:0] ? myVec_72 : _GEN_15601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15603 = 7'h49 == _myNewVec_7_T_3[6:0] ? myVec_73 : _GEN_15602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15604 = 7'h4a == _myNewVec_7_T_3[6:0] ? myVec_74 : _GEN_15603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15605 = 7'h4b == _myNewVec_7_T_3[6:0] ? myVec_75 : _GEN_15604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15606 = 7'h4c == _myNewVec_7_T_3[6:0] ? myVec_76 : _GEN_15605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15607 = 7'h4d == _myNewVec_7_T_3[6:0] ? myVec_77 : _GEN_15606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15608 = 7'h4e == _myNewVec_7_T_3[6:0] ? myVec_78 : _GEN_15607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15609 = 7'h4f == _myNewVec_7_T_3[6:0] ? myVec_79 : _GEN_15608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15610 = 7'h50 == _myNewVec_7_T_3[6:0] ? myVec_80 : _GEN_15609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15611 = 7'h51 == _myNewVec_7_T_3[6:0] ? myVec_81 : _GEN_15610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15612 = 7'h52 == _myNewVec_7_T_3[6:0] ? myVec_82 : _GEN_15611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15613 = 7'h53 == _myNewVec_7_T_3[6:0] ? myVec_83 : _GEN_15612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15614 = 7'h54 == _myNewVec_7_T_3[6:0] ? myVec_84 : _GEN_15613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15615 = 7'h55 == _myNewVec_7_T_3[6:0] ? myVec_85 : _GEN_15614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15616 = 7'h56 == _myNewVec_7_T_3[6:0] ? myVec_86 : _GEN_15615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15617 = 7'h57 == _myNewVec_7_T_3[6:0] ? myVec_87 : _GEN_15616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15618 = 7'h58 == _myNewVec_7_T_3[6:0] ? myVec_88 : _GEN_15617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15619 = 7'h59 == _myNewVec_7_T_3[6:0] ? myVec_89 : _GEN_15618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15620 = 7'h5a == _myNewVec_7_T_3[6:0] ? myVec_90 : _GEN_15619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15621 = 7'h5b == _myNewVec_7_T_3[6:0] ? myVec_91 : _GEN_15620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15622 = 7'h5c == _myNewVec_7_T_3[6:0] ? myVec_92 : _GEN_15621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15623 = 7'h5d == _myNewVec_7_T_3[6:0] ? myVec_93 : _GEN_15622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15624 = 7'h5e == _myNewVec_7_T_3[6:0] ? myVec_94 : _GEN_15623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15625 = 7'h5f == _myNewVec_7_T_3[6:0] ? myVec_95 : _GEN_15624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15626 = 7'h60 == _myNewVec_7_T_3[6:0] ? myVec_96 : _GEN_15625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15627 = 7'h61 == _myNewVec_7_T_3[6:0] ? myVec_97 : _GEN_15626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15628 = 7'h62 == _myNewVec_7_T_3[6:0] ? myVec_98 : _GEN_15627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15629 = 7'h63 == _myNewVec_7_T_3[6:0] ? myVec_99 : _GEN_15628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15630 = 7'h64 == _myNewVec_7_T_3[6:0] ? myVec_100 : _GEN_15629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15631 = 7'h65 == _myNewVec_7_T_3[6:0] ? myVec_101 : _GEN_15630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15632 = 7'h66 == _myNewVec_7_T_3[6:0] ? myVec_102 : _GEN_15631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15633 = 7'h67 == _myNewVec_7_T_3[6:0] ? myVec_103 : _GEN_15632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15634 = 7'h68 == _myNewVec_7_T_3[6:0] ? myVec_104 : _GEN_15633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15635 = 7'h69 == _myNewVec_7_T_3[6:0] ? myVec_105 : _GEN_15634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15636 = 7'h6a == _myNewVec_7_T_3[6:0] ? myVec_106 : _GEN_15635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15637 = 7'h6b == _myNewVec_7_T_3[6:0] ? myVec_107 : _GEN_15636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15638 = 7'h6c == _myNewVec_7_T_3[6:0] ? myVec_108 : _GEN_15637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15639 = 7'h6d == _myNewVec_7_T_3[6:0] ? myVec_109 : _GEN_15638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15640 = 7'h6e == _myNewVec_7_T_3[6:0] ? myVec_110 : _GEN_15639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15641 = 7'h6f == _myNewVec_7_T_3[6:0] ? myVec_111 : _GEN_15640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15642 = 7'h70 == _myNewVec_7_T_3[6:0] ? myVec_112 : _GEN_15641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15643 = 7'h71 == _myNewVec_7_T_3[6:0] ? myVec_113 : _GEN_15642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15644 = 7'h72 == _myNewVec_7_T_3[6:0] ? myVec_114 : _GEN_15643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15645 = 7'h73 == _myNewVec_7_T_3[6:0] ? myVec_115 : _GEN_15644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15646 = 7'h74 == _myNewVec_7_T_3[6:0] ? myVec_116 : _GEN_15645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15647 = 7'h75 == _myNewVec_7_T_3[6:0] ? myVec_117 : _GEN_15646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15648 = 7'h76 == _myNewVec_7_T_3[6:0] ? myVec_118 : _GEN_15647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15649 = 7'h77 == _myNewVec_7_T_3[6:0] ? myVec_119 : _GEN_15648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15650 = 7'h78 == _myNewVec_7_T_3[6:0] ? myVec_120 : _GEN_15649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15651 = 7'h79 == _myNewVec_7_T_3[6:0] ? myVec_121 : _GEN_15650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15652 = 7'h7a == _myNewVec_7_T_3[6:0] ? myVec_122 : _GEN_15651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15653 = 7'h7b == _myNewVec_7_T_3[6:0] ? myVec_123 : _GEN_15652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15654 = 7'h7c == _myNewVec_7_T_3[6:0] ? myVec_124 : _GEN_15653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15655 = 7'h7d == _myNewVec_7_T_3[6:0] ? myVec_125 : _GEN_15654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15656 = 7'h7e == _myNewVec_7_T_3[6:0] ? myVec_126 : _GEN_15655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_7 = 7'h7f == _myNewVec_7_T_3[6:0] ? myVec_127 : _GEN_15656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_6_T_3 = _myNewVec_127_T_1 + 16'h79; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_15659 = 7'h1 == _myNewVec_6_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15660 = 7'h2 == _myNewVec_6_T_3[6:0] ? myVec_2 : _GEN_15659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15661 = 7'h3 == _myNewVec_6_T_3[6:0] ? myVec_3 : _GEN_15660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15662 = 7'h4 == _myNewVec_6_T_3[6:0] ? myVec_4 : _GEN_15661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15663 = 7'h5 == _myNewVec_6_T_3[6:0] ? myVec_5 : _GEN_15662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15664 = 7'h6 == _myNewVec_6_T_3[6:0] ? myVec_6 : _GEN_15663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15665 = 7'h7 == _myNewVec_6_T_3[6:0] ? myVec_7 : _GEN_15664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15666 = 7'h8 == _myNewVec_6_T_3[6:0] ? myVec_8 : _GEN_15665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15667 = 7'h9 == _myNewVec_6_T_3[6:0] ? myVec_9 : _GEN_15666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15668 = 7'ha == _myNewVec_6_T_3[6:0] ? myVec_10 : _GEN_15667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15669 = 7'hb == _myNewVec_6_T_3[6:0] ? myVec_11 : _GEN_15668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15670 = 7'hc == _myNewVec_6_T_3[6:0] ? myVec_12 : _GEN_15669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15671 = 7'hd == _myNewVec_6_T_3[6:0] ? myVec_13 : _GEN_15670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15672 = 7'he == _myNewVec_6_T_3[6:0] ? myVec_14 : _GEN_15671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15673 = 7'hf == _myNewVec_6_T_3[6:0] ? myVec_15 : _GEN_15672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15674 = 7'h10 == _myNewVec_6_T_3[6:0] ? myVec_16 : _GEN_15673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15675 = 7'h11 == _myNewVec_6_T_3[6:0] ? myVec_17 : _GEN_15674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15676 = 7'h12 == _myNewVec_6_T_3[6:0] ? myVec_18 : _GEN_15675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15677 = 7'h13 == _myNewVec_6_T_3[6:0] ? myVec_19 : _GEN_15676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15678 = 7'h14 == _myNewVec_6_T_3[6:0] ? myVec_20 : _GEN_15677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15679 = 7'h15 == _myNewVec_6_T_3[6:0] ? myVec_21 : _GEN_15678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15680 = 7'h16 == _myNewVec_6_T_3[6:0] ? myVec_22 : _GEN_15679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15681 = 7'h17 == _myNewVec_6_T_3[6:0] ? myVec_23 : _GEN_15680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15682 = 7'h18 == _myNewVec_6_T_3[6:0] ? myVec_24 : _GEN_15681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15683 = 7'h19 == _myNewVec_6_T_3[6:0] ? myVec_25 : _GEN_15682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15684 = 7'h1a == _myNewVec_6_T_3[6:0] ? myVec_26 : _GEN_15683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15685 = 7'h1b == _myNewVec_6_T_3[6:0] ? myVec_27 : _GEN_15684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15686 = 7'h1c == _myNewVec_6_T_3[6:0] ? myVec_28 : _GEN_15685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15687 = 7'h1d == _myNewVec_6_T_3[6:0] ? myVec_29 : _GEN_15686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15688 = 7'h1e == _myNewVec_6_T_3[6:0] ? myVec_30 : _GEN_15687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15689 = 7'h1f == _myNewVec_6_T_3[6:0] ? myVec_31 : _GEN_15688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15690 = 7'h20 == _myNewVec_6_T_3[6:0] ? myVec_32 : _GEN_15689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15691 = 7'h21 == _myNewVec_6_T_3[6:0] ? myVec_33 : _GEN_15690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15692 = 7'h22 == _myNewVec_6_T_3[6:0] ? myVec_34 : _GEN_15691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15693 = 7'h23 == _myNewVec_6_T_3[6:0] ? myVec_35 : _GEN_15692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15694 = 7'h24 == _myNewVec_6_T_3[6:0] ? myVec_36 : _GEN_15693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15695 = 7'h25 == _myNewVec_6_T_3[6:0] ? myVec_37 : _GEN_15694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15696 = 7'h26 == _myNewVec_6_T_3[6:0] ? myVec_38 : _GEN_15695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15697 = 7'h27 == _myNewVec_6_T_3[6:0] ? myVec_39 : _GEN_15696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15698 = 7'h28 == _myNewVec_6_T_3[6:0] ? myVec_40 : _GEN_15697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15699 = 7'h29 == _myNewVec_6_T_3[6:0] ? myVec_41 : _GEN_15698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15700 = 7'h2a == _myNewVec_6_T_3[6:0] ? myVec_42 : _GEN_15699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15701 = 7'h2b == _myNewVec_6_T_3[6:0] ? myVec_43 : _GEN_15700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15702 = 7'h2c == _myNewVec_6_T_3[6:0] ? myVec_44 : _GEN_15701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15703 = 7'h2d == _myNewVec_6_T_3[6:0] ? myVec_45 : _GEN_15702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15704 = 7'h2e == _myNewVec_6_T_3[6:0] ? myVec_46 : _GEN_15703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15705 = 7'h2f == _myNewVec_6_T_3[6:0] ? myVec_47 : _GEN_15704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15706 = 7'h30 == _myNewVec_6_T_3[6:0] ? myVec_48 : _GEN_15705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15707 = 7'h31 == _myNewVec_6_T_3[6:0] ? myVec_49 : _GEN_15706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15708 = 7'h32 == _myNewVec_6_T_3[6:0] ? myVec_50 : _GEN_15707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15709 = 7'h33 == _myNewVec_6_T_3[6:0] ? myVec_51 : _GEN_15708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15710 = 7'h34 == _myNewVec_6_T_3[6:0] ? myVec_52 : _GEN_15709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15711 = 7'h35 == _myNewVec_6_T_3[6:0] ? myVec_53 : _GEN_15710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15712 = 7'h36 == _myNewVec_6_T_3[6:0] ? myVec_54 : _GEN_15711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15713 = 7'h37 == _myNewVec_6_T_3[6:0] ? myVec_55 : _GEN_15712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15714 = 7'h38 == _myNewVec_6_T_3[6:0] ? myVec_56 : _GEN_15713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15715 = 7'h39 == _myNewVec_6_T_3[6:0] ? myVec_57 : _GEN_15714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15716 = 7'h3a == _myNewVec_6_T_3[6:0] ? myVec_58 : _GEN_15715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15717 = 7'h3b == _myNewVec_6_T_3[6:0] ? myVec_59 : _GEN_15716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15718 = 7'h3c == _myNewVec_6_T_3[6:0] ? myVec_60 : _GEN_15717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15719 = 7'h3d == _myNewVec_6_T_3[6:0] ? myVec_61 : _GEN_15718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15720 = 7'h3e == _myNewVec_6_T_3[6:0] ? myVec_62 : _GEN_15719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15721 = 7'h3f == _myNewVec_6_T_3[6:0] ? myVec_63 : _GEN_15720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15722 = 7'h40 == _myNewVec_6_T_3[6:0] ? myVec_64 : _GEN_15721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15723 = 7'h41 == _myNewVec_6_T_3[6:0] ? myVec_65 : _GEN_15722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15724 = 7'h42 == _myNewVec_6_T_3[6:0] ? myVec_66 : _GEN_15723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15725 = 7'h43 == _myNewVec_6_T_3[6:0] ? myVec_67 : _GEN_15724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15726 = 7'h44 == _myNewVec_6_T_3[6:0] ? myVec_68 : _GEN_15725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15727 = 7'h45 == _myNewVec_6_T_3[6:0] ? myVec_69 : _GEN_15726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15728 = 7'h46 == _myNewVec_6_T_3[6:0] ? myVec_70 : _GEN_15727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15729 = 7'h47 == _myNewVec_6_T_3[6:0] ? myVec_71 : _GEN_15728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15730 = 7'h48 == _myNewVec_6_T_3[6:0] ? myVec_72 : _GEN_15729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15731 = 7'h49 == _myNewVec_6_T_3[6:0] ? myVec_73 : _GEN_15730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15732 = 7'h4a == _myNewVec_6_T_3[6:0] ? myVec_74 : _GEN_15731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15733 = 7'h4b == _myNewVec_6_T_3[6:0] ? myVec_75 : _GEN_15732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15734 = 7'h4c == _myNewVec_6_T_3[6:0] ? myVec_76 : _GEN_15733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15735 = 7'h4d == _myNewVec_6_T_3[6:0] ? myVec_77 : _GEN_15734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15736 = 7'h4e == _myNewVec_6_T_3[6:0] ? myVec_78 : _GEN_15735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15737 = 7'h4f == _myNewVec_6_T_3[6:0] ? myVec_79 : _GEN_15736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15738 = 7'h50 == _myNewVec_6_T_3[6:0] ? myVec_80 : _GEN_15737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15739 = 7'h51 == _myNewVec_6_T_3[6:0] ? myVec_81 : _GEN_15738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15740 = 7'h52 == _myNewVec_6_T_3[6:0] ? myVec_82 : _GEN_15739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15741 = 7'h53 == _myNewVec_6_T_3[6:0] ? myVec_83 : _GEN_15740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15742 = 7'h54 == _myNewVec_6_T_3[6:0] ? myVec_84 : _GEN_15741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15743 = 7'h55 == _myNewVec_6_T_3[6:0] ? myVec_85 : _GEN_15742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15744 = 7'h56 == _myNewVec_6_T_3[6:0] ? myVec_86 : _GEN_15743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15745 = 7'h57 == _myNewVec_6_T_3[6:0] ? myVec_87 : _GEN_15744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15746 = 7'h58 == _myNewVec_6_T_3[6:0] ? myVec_88 : _GEN_15745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15747 = 7'h59 == _myNewVec_6_T_3[6:0] ? myVec_89 : _GEN_15746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15748 = 7'h5a == _myNewVec_6_T_3[6:0] ? myVec_90 : _GEN_15747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15749 = 7'h5b == _myNewVec_6_T_3[6:0] ? myVec_91 : _GEN_15748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15750 = 7'h5c == _myNewVec_6_T_3[6:0] ? myVec_92 : _GEN_15749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15751 = 7'h5d == _myNewVec_6_T_3[6:0] ? myVec_93 : _GEN_15750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15752 = 7'h5e == _myNewVec_6_T_3[6:0] ? myVec_94 : _GEN_15751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15753 = 7'h5f == _myNewVec_6_T_3[6:0] ? myVec_95 : _GEN_15752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15754 = 7'h60 == _myNewVec_6_T_3[6:0] ? myVec_96 : _GEN_15753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15755 = 7'h61 == _myNewVec_6_T_3[6:0] ? myVec_97 : _GEN_15754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15756 = 7'h62 == _myNewVec_6_T_3[6:0] ? myVec_98 : _GEN_15755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15757 = 7'h63 == _myNewVec_6_T_3[6:0] ? myVec_99 : _GEN_15756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15758 = 7'h64 == _myNewVec_6_T_3[6:0] ? myVec_100 : _GEN_15757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15759 = 7'h65 == _myNewVec_6_T_3[6:0] ? myVec_101 : _GEN_15758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15760 = 7'h66 == _myNewVec_6_T_3[6:0] ? myVec_102 : _GEN_15759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15761 = 7'h67 == _myNewVec_6_T_3[6:0] ? myVec_103 : _GEN_15760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15762 = 7'h68 == _myNewVec_6_T_3[6:0] ? myVec_104 : _GEN_15761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15763 = 7'h69 == _myNewVec_6_T_3[6:0] ? myVec_105 : _GEN_15762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15764 = 7'h6a == _myNewVec_6_T_3[6:0] ? myVec_106 : _GEN_15763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15765 = 7'h6b == _myNewVec_6_T_3[6:0] ? myVec_107 : _GEN_15764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15766 = 7'h6c == _myNewVec_6_T_3[6:0] ? myVec_108 : _GEN_15765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15767 = 7'h6d == _myNewVec_6_T_3[6:0] ? myVec_109 : _GEN_15766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15768 = 7'h6e == _myNewVec_6_T_3[6:0] ? myVec_110 : _GEN_15767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15769 = 7'h6f == _myNewVec_6_T_3[6:0] ? myVec_111 : _GEN_15768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15770 = 7'h70 == _myNewVec_6_T_3[6:0] ? myVec_112 : _GEN_15769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15771 = 7'h71 == _myNewVec_6_T_3[6:0] ? myVec_113 : _GEN_15770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15772 = 7'h72 == _myNewVec_6_T_3[6:0] ? myVec_114 : _GEN_15771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15773 = 7'h73 == _myNewVec_6_T_3[6:0] ? myVec_115 : _GEN_15772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15774 = 7'h74 == _myNewVec_6_T_3[6:0] ? myVec_116 : _GEN_15773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15775 = 7'h75 == _myNewVec_6_T_3[6:0] ? myVec_117 : _GEN_15774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15776 = 7'h76 == _myNewVec_6_T_3[6:0] ? myVec_118 : _GEN_15775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15777 = 7'h77 == _myNewVec_6_T_3[6:0] ? myVec_119 : _GEN_15776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15778 = 7'h78 == _myNewVec_6_T_3[6:0] ? myVec_120 : _GEN_15777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15779 = 7'h79 == _myNewVec_6_T_3[6:0] ? myVec_121 : _GEN_15778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15780 = 7'h7a == _myNewVec_6_T_3[6:0] ? myVec_122 : _GEN_15779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15781 = 7'h7b == _myNewVec_6_T_3[6:0] ? myVec_123 : _GEN_15780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15782 = 7'h7c == _myNewVec_6_T_3[6:0] ? myVec_124 : _GEN_15781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15783 = 7'h7d == _myNewVec_6_T_3[6:0] ? myVec_125 : _GEN_15782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15784 = 7'h7e == _myNewVec_6_T_3[6:0] ? myVec_126 : _GEN_15783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_6 = 7'h7f == _myNewVec_6_T_3[6:0] ? myVec_127 : _GEN_15784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_5_T_3 = _myNewVec_127_T_1 + 16'h7a; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_15787 = 7'h1 == _myNewVec_5_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15788 = 7'h2 == _myNewVec_5_T_3[6:0] ? myVec_2 : _GEN_15787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15789 = 7'h3 == _myNewVec_5_T_3[6:0] ? myVec_3 : _GEN_15788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15790 = 7'h4 == _myNewVec_5_T_3[6:0] ? myVec_4 : _GEN_15789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15791 = 7'h5 == _myNewVec_5_T_3[6:0] ? myVec_5 : _GEN_15790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15792 = 7'h6 == _myNewVec_5_T_3[6:0] ? myVec_6 : _GEN_15791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15793 = 7'h7 == _myNewVec_5_T_3[6:0] ? myVec_7 : _GEN_15792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15794 = 7'h8 == _myNewVec_5_T_3[6:0] ? myVec_8 : _GEN_15793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15795 = 7'h9 == _myNewVec_5_T_3[6:0] ? myVec_9 : _GEN_15794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15796 = 7'ha == _myNewVec_5_T_3[6:0] ? myVec_10 : _GEN_15795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15797 = 7'hb == _myNewVec_5_T_3[6:0] ? myVec_11 : _GEN_15796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15798 = 7'hc == _myNewVec_5_T_3[6:0] ? myVec_12 : _GEN_15797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15799 = 7'hd == _myNewVec_5_T_3[6:0] ? myVec_13 : _GEN_15798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15800 = 7'he == _myNewVec_5_T_3[6:0] ? myVec_14 : _GEN_15799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15801 = 7'hf == _myNewVec_5_T_3[6:0] ? myVec_15 : _GEN_15800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15802 = 7'h10 == _myNewVec_5_T_3[6:0] ? myVec_16 : _GEN_15801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15803 = 7'h11 == _myNewVec_5_T_3[6:0] ? myVec_17 : _GEN_15802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15804 = 7'h12 == _myNewVec_5_T_3[6:0] ? myVec_18 : _GEN_15803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15805 = 7'h13 == _myNewVec_5_T_3[6:0] ? myVec_19 : _GEN_15804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15806 = 7'h14 == _myNewVec_5_T_3[6:0] ? myVec_20 : _GEN_15805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15807 = 7'h15 == _myNewVec_5_T_3[6:0] ? myVec_21 : _GEN_15806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15808 = 7'h16 == _myNewVec_5_T_3[6:0] ? myVec_22 : _GEN_15807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15809 = 7'h17 == _myNewVec_5_T_3[6:0] ? myVec_23 : _GEN_15808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15810 = 7'h18 == _myNewVec_5_T_3[6:0] ? myVec_24 : _GEN_15809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15811 = 7'h19 == _myNewVec_5_T_3[6:0] ? myVec_25 : _GEN_15810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15812 = 7'h1a == _myNewVec_5_T_3[6:0] ? myVec_26 : _GEN_15811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15813 = 7'h1b == _myNewVec_5_T_3[6:0] ? myVec_27 : _GEN_15812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15814 = 7'h1c == _myNewVec_5_T_3[6:0] ? myVec_28 : _GEN_15813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15815 = 7'h1d == _myNewVec_5_T_3[6:0] ? myVec_29 : _GEN_15814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15816 = 7'h1e == _myNewVec_5_T_3[6:0] ? myVec_30 : _GEN_15815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15817 = 7'h1f == _myNewVec_5_T_3[6:0] ? myVec_31 : _GEN_15816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15818 = 7'h20 == _myNewVec_5_T_3[6:0] ? myVec_32 : _GEN_15817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15819 = 7'h21 == _myNewVec_5_T_3[6:0] ? myVec_33 : _GEN_15818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15820 = 7'h22 == _myNewVec_5_T_3[6:0] ? myVec_34 : _GEN_15819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15821 = 7'h23 == _myNewVec_5_T_3[6:0] ? myVec_35 : _GEN_15820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15822 = 7'h24 == _myNewVec_5_T_3[6:0] ? myVec_36 : _GEN_15821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15823 = 7'h25 == _myNewVec_5_T_3[6:0] ? myVec_37 : _GEN_15822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15824 = 7'h26 == _myNewVec_5_T_3[6:0] ? myVec_38 : _GEN_15823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15825 = 7'h27 == _myNewVec_5_T_3[6:0] ? myVec_39 : _GEN_15824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15826 = 7'h28 == _myNewVec_5_T_3[6:0] ? myVec_40 : _GEN_15825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15827 = 7'h29 == _myNewVec_5_T_3[6:0] ? myVec_41 : _GEN_15826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15828 = 7'h2a == _myNewVec_5_T_3[6:0] ? myVec_42 : _GEN_15827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15829 = 7'h2b == _myNewVec_5_T_3[6:0] ? myVec_43 : _GEN_15828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15830 = 7'h2c == _myNewVec_5_T_3[6:0] ? myVec_44 : _GEN_15829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15831 = 7'h2d == _myNewVec_5_T_3[6:0] ? myVec_45 : _GEN_15830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15832 = 7'h2e == _myNewVec_5_T_3[6:0] ? myVec_46 : _GEN_15831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15833 = 7'h2f == _myNewVec_5_T_3[6:0] ? myVec_47 : _GEN_15832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15834 = 7'h30 == _myNewVec_5_T_3[6:0] ? myVec_48 : _GEN_15833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15835 = 7'h31 == _myNewVec_5_T_3[6:0] ? myVec_49 : _GEN_15834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15836 = 7'h32 == _myNewVec_5_T_3[6:0] ? myVec_50 : _GEN_15835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15837 = 7'h33 == _myNewVec_5_T_3[6:0] ? myVec_51 : _GEN_15836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15838 = 7'h34 == _myNewVec_5_T_3[6:0] ? myVec_52 : _GEN_15837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15839 = 7'h35 == _myNewVec_5_T_3[6:0] ? myVec_53 : _GEN_15838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15840 = 7'h36 == _myNewVec_5_T_3[6:0] ? myVec_54 : _GEN_15839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15841 = 7'h37 == _myNewVec_5_T_3[6:0] ? myVec_55 : _GEN_15840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15842 = 7'h38 == _myNewVec_5_T_3[6:0] ? myVec_56 : _GEN_15841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15843 = 7'h39 == _myNewVec_5_T_3[6:0] ? myVec_57 : _GEN_15842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15844 = 7'h3a == _myNewVec_5_T_3[6:0] ? myVec_58 : _GEN_15843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15845 = 7'h3b == _myNewVec_5_T_3[6:0] ? myVec_59 : _GEN_15844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15846 = 7'h3c == _myNewVec_5_T_3[6:0] ? myVec_60 : _GEN_15845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15847 = 7'h3d == _myNewVec_5_T_3[6:0] ? myVec_61 : _GEN_15846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15848 = 7'h3e == _myNewVec_5_T_3[6:0] ? myVec_62 : _GEN_15847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15849 = 7'h3f == _myNewVec_5_T_3[6:0] ? myVec_63 : _GEN_15848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15850 = 7'h40 == _myNewVec_5_T_3[6:0] ? myVec_64 : _GEN_15849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15851 = 7'h41 == _myNewVec_5_T_3[6:0] ? myVec_65 : _GEN_15850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15852 = 7'h42 == _myNewVec_5_T_3[6:0] ? myVec_66 : _GEN_15851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15853 = 7'h43 == _myNewVec_5_T_3[6:0] ? myVec_67 : _GEN_15852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15854 = 7'h44 == _myNewVec_5_T_3[6:0] ? myVec_68 : _GEN_15853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15855 = 7'h45 == _myNewVec_5_T_3[6:0] ? myVec_69 : _GEN_15854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15856 = 7'h46 == _myNewVec_5_T_3[6:0] ? myVec_70 : _GEN_15855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15857 = 7'h47 == _myNewVec_5_T_3[6:0] ? myVec_71 : _GEN_15856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15858 = 7'h48 == _myNewVec_5_T_3[6:0] ? myVec_72 : _GEN_15857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15859 = 7'h49 == _myNewVec_5_T_3[6:0] ? myVec_73 : _GEN_15858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15860 = 7'h4a == _myNewVec_5_T_3[6:0] ? myVec_74 : _GEN_15859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15861 = 7'h4b == _myNewVec_5_T_3[6:0] ? myVec_75 : _GEN_15860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15862 = 7'h4c == _myNewVec_5_T_3[6:0] ? myVec_76 : _GEN_15861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15863 = 7'h4d == _myNewVec_5_T_3[6:0] ? myVec_77 : _GEN_15862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15864 = 7'h4e == _myNewVec_5_T_3[6:0] ? myVec_78 : _GEN_15863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15865 = 7'h4f == _myNewVec_5_T_3[6:0] ? myVec_79 : _GEN_15864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15866 = 7'h50 == _myNewVec_5_T_3[6:0] ? myVec_80 : _GEN_15865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15867 = 7'h51 == _myNewVec_5_T_3[6:0] ? myVec_81 : _GEN_15866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15868 = 7'h52 == _myNewVec_5_T_3[6:0] ? myVec_82 : _GEN_15867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15869 = 7'h53 == _myNewVec_5_T_3[6:0] ? myVec_83 : _GEN_15868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15870 = 7'h54 == _myNewVec_5_T_3[6:0] ? myVec_84 : _GEN_15869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15871 = 7'h55 == _myNewVec_5_T_3[6:0] ? myVec_85 : _GEN_15870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15872 = 7'h56 == _myNewVec_5_T_3[6:0] ? myVec_86 : _GEN_15871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15873 = 7'h57 == _myNewVec_5_T_3[6:0] ? myVec_87 : _GEN_15872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15874 = 7'h58 == _myNewVec_5_T_3[6:0] ? myVec_88 : _GEN_15873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15875 = 7'h59 == _myNewVec_5_T_3[6:0] ? myVec_89 : _GEN_15874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15876 = 7'h5a == _myNewVec_5_T_3[6:0] ? myVec_90 : _GEN_15875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15877 = 7'h5b == _myNewVec_5_T_3[6:0] ? myVec_91 : _GEN_15876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15878 = 7'h5c == _myNewVec_5_T_3[6:0] ? myVec_92 : _GEN_15877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15879 = 7'h5d == _myNewVec_5_T_3[6:0] ? myVec_93 : _GEN_15878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15880 = 7'h5e == _myNewVec_5_T_3[6:0] ? myVec_94 : _GEN_15879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15881 = 7'h5f == _myNewVec_5_T_3[6:0] ? myVec_95 : _GEN_15880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15882 = 7'h60 == _myNewVec_5_T_3[6:0] ? myVec_96 : _GEN_15881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15883 = 7'h61 == _myNewVec_5_T_3[6:0] ? myVec_97 : _GEN_15882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15884 = 7'h62 == _myNewVec_5_T_3[6:0] ? myVec_98 : _GEN_15883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15885 = 7'h63 == _myNewVec_5_T_3[6:0] ? myVec_99 : _GEN_15884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15886 = 7'h64 == _myNewVec_5_T_3[6:0] ? myVec_100 : _GEN_15885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15887 = 7'h65 == _myNewVec_5_T_3[6:0] ? myVec_101 : _GEN_15886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15888 = 7'h66 == _myNewVec_5_T_3[6:0] ? myVec_102 : _GEN_15887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15889 = 7'h67 == _myNewVec_5_T_3[6:0] ? myVec_103 : _GEN_15888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15890 = 7'h68 == _myNewVec_5_T_3[6:0] ? myVec_104 : _GEN_15889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15891 = 7'h69 == _myNewVec_5_T_3[6:0] ? myVec_105 : _GEN_15890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15892 = 7'h6a == _myNewVec_5_T_3[6:0] ? myVec_106 : _GEN_15891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15893 = 7'h6b == _myNewVec_5_T_3[6:0] ? myVec_107 : _GEN_15892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15894 = 7'h6c == _myNewVec_5_T_3[6:0] ? myVec_108 : _GEN_15893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15895 = 7'h6d == _myNewVec_5_T_3[6:0] ? myVec_109 : _GEN_15894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15896 = 7'h6e == _myNewVec_5_T_3[6:0] ? myVec_110 : _GEN_15895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15897 = 7'h6f == _myNewVec_5_T_3[6:0] ? myVec_111 : _GEN_15896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15898 = 7'h70 == _myNewVec_5_T_3[6:0] ? myVec_112 : _GEN_15897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15899 = 7'h71 == _myNewVec_5_T_3[6:0] ? myVec_113 : _GEN_15898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15900 = 7'h72 == _myNewVec_5_T_3[6:0] ? myVec_114 : _GEN_15899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15901 = 7'h73 == _myNewVec_5_T_3[6:0] ? myVec_115 : _GEN_15900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15902 = 7'h74 == _myNewVec_5_T_3[6:0] ? myVec_116 : _GEN_15901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15903 = 7'h75 == _myNewVec_5_T_3[6:0] ? myVec_117 : _GEN_15902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15904 = 7'h76 == _myNewVec_5_T_3[6:0] ? myVec_118 : _GEN_15903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15905 = 7'h77 == _myNewVec_5_T_3[6:0] ? myVec_119 : _GEN_15904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15906 = 7'h78 == _myNewVec_5_T_3[6:0] ? myVec_120 : _GEN_15905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15907 = 7'h79 == _myNewVec_5_T_3[6:0] ? myVec_121 : _GEN_15906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15908 = 7'h7a == _myNewVec_5_T_3[6:0] ? myVec_122 : _GEN_15907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15909 = 7'h7b == _myNewVec_5_T_3[6:0] ? myVec_123 : _GEN_15908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15910 = 7'h7c == _myNewVec_5_T_3[6:0] ? myVec_124 : _GEN_15909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15911 = 7'h7d == _myNewVec_5_T_3[6:0] ? myVec_125 : _GEN_15910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15912 = 7'h7e == _myNewVec_5_T_3[6:0] ? myVec_126 : _GEN_15911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_5 = 7'h7f == _myNewVec_5_T_3[6:0] ? myVec_127 : _GEN_15912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_4_T_3 = _myNewVec_127_T_1 + 16'h7b; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_15915 = 7'h1 == _myNewVec_4_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15916 = 7'h2 == _myNewVec_4_T_3[6:0] ? myVec_2 : _GEN_15915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15917 = 7'h3 == _myNewVec_4_T_3[6:0] ? myVec_3 : _GEN_15916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15918 = 7'h4 == _myNewVec_4_T_3[6:0] ? myVec_4 : _GEN_15917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15919 = 7'h5 == _myNewVec_4_T_3[6:0] ? myVec_5 : _GEN_15918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15920 = 7'h6 == _myNewVec_4_T_3[6:0] ? myVec_6 : _GEN_15919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15921 = 7'h7 == _myNewVec_4_T_3[6:0] ? myVec_7 : _GEN_15920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15922 = 7'h8 == _myNewVec_4_T_3[6:0] ? myVec_8 : _GEN_15921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15923 = 7'h9 == _myNewVec_4_T_3[6:0] ? myVec_9 : _GEN_15922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15924 = 7'ha == _myNewVec_4_T_3[6:0] ? myVec_10 : _GEN_15923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15925 = 7'hb == _myNewVec_4_T_3[6:0] ? myVec_11 : _GEN_15924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15926 = 7'hc == _myNewVec_4_T_3[6:0] ? myVec_12 : _GEN_15925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15927 = 7'hd == _myNewVec_4_T_3[6:0] ? myVec_13 : _GEN_15926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15928 = 7'he == _myNewVec_4_T_3[6:0] ? myVec_14 : _GEN_15927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15929 = 7'hf == _myNewVec_4_T_3[6:0] ? myVec_15 : _GEN_15928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15930 = 7'h10 == _myNewVec_4_T_3[6:0] ? myVec_16 : _GEN_15929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15931 = 7'h11 == _myNewVec_4_T_3[6:0] ? myVec_17 : _GEN_15930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15932 = 7'h12 == _myNewVec_4_T_3[6:0] ? myVec_18 : _GEN_15931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15933 = 7'h13 == _myNewVec_4_T_3[6:0] ? myVec_19 : _GEN_15932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15934 = 7'h14 == _myNewVec_4_T_3[6:0] ? myVec_20 : _GEN_15933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15935 = 7'h15 == _myNewVec_4_T_3[6:0] ? myVec_21 : _GEN_15934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15936 = 7'h16 == _myNewVec_4_T_3[6:0] ? myVec_22 : _GEN_15935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15937 = 7'h17 == _myNewVec_4_T_3[6:0] ? myVec_23 : _GEN_15936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15938 = 7'h18 == _myNewVec_4_T_3[6:0] ? myVec_24 : _GEN_15937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15939 = 7'h19 == _myNewVec_4_T_3[6:0] ? myVec_25 : _GEN_15938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15940 = 7'h1a == _myNewVec_4_T_3[6:0] ? myVec_26 : _GEN_15939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15941 = 7'h1b == _myNewVec_4_T_3[6:0] ? myVec_27 : _GEN_15940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15942 = 7'h1c == _myNewVec_4_T_3[6:0] ? myVec_28 : _GEN_15941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15943 = 7'h1d == _myNewVec_4_T_3[6:0] ? myVec_29 : _GEN_15942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15944 = 7'h1e == _myNewVec_4_T_3[6:0] ? myVec_30 : _GEN_15943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15945 = 7'h1f == _myNewVec_4_T_3[6:0] ? myVec_31 : _GEN_15944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15946 = 7'h20 == _myNewVec_4_T_3[6:0] ? myVec_32 : _GEN_15945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15947 = 7'h21 == _myNewVec_4_T_3[6:0] ? myVec_33 : _GEN_15946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15948 = 7'h22 == _myNewVec_4_T_3[6:0] ? myVec_34 : _GEN_15947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15949 = 7'h23 == _myNewVec_4_T_3[6:0] ? myVec_35 : _GEN_15948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15950 = 7'h24 == _myNewVec_4_T_3[6:0] ? myVec_36 : _GEN_15949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15951 = 7'h25 == _myNewVec_4_T_3[6:0] ? myVec_37 : _GEN_15950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15952 = 7'h26 == _myNewVec_4_T_3[6:0] ? myVec_38 : _GEN_15951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15953 = 7'h27 == _myNewVec_4_T_3[6:0] ? myVec_39 : _GEN_15952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15954 = 7'h28 == _myNewVec_4_T_3[6:0] ? myVec_40 : _GEN_15953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15955 = 7'h29 == _myNewVec_4_T_3[6:0] ? myVec_41 : _GEN_15954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15956 = 7'h2a == _myNewVec_4_T_3[6:0] ? myVec_42 : _GEN_15955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15957 = 7'h2b == _myNewVec_4_T_3[6:0] ? myVec_43 : _GEN_15956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15958 = 7'h2c == _myNewVec_4_T_3[6:0] ? myVec_44 : _GEN_15957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15959 = 7'h2d == _myNewVec_4_T_3[6:0] ? myVec_45 : _GEN_15958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15960 = 7'h2e == _myNewVec_4_T_3[6:0] ? myVec_46 : _GEN_15959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15961 = 7'h2f == _myNewVec_4_T_3[6:0] ? myVec_47 : _GEN_15960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15962 = 7'h30 == _myNewVec_4_T_3[6:0] ? myVec_48 : _GEN_15961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15963 = 7'h31 == _myNewVec_4_T_3[6:0] ? myVec_49 : _GEN_15962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15964 = 7'h32 == _myNewVec_4_T_3[6:0] ? myVec_50 : _GEN_15963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15965 = 7'h33 == _myNewVec_4_T_3[6:0] ? myVec_51 : _GEN_15964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15966 = 7'h34 == _myNewVec_4_T_3[6:0] ? myVec_52 : _GEN_15965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15967 = 7'h35 == _myNewVec_4_T_3[6:0] ? myVec_53 : _GEN_15966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15968 = 7'h36 == _myNewVec_4_T_3[6:0] ? myVec_54 : _GEN_15967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15969 = 7'h37 == _myNewVec_4_T_3[6:0] ? myVec_55 : _GEN_15968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15970 = 7'h38 == _myNewVec_4_T_3[6:0] ? myVec_56 : _GEN_15969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15971 = 7'h39 == _myNewVec_4_T_3[6:0] ? myVec_57 : _GEN_15970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15972 = 7'h3a == _myNewVec_4_T_3[6:0] ? myVec_58 : _GEN_15971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15973 = 7'h3b == _myNewVec_4_T_3[6:0] ? myVec_59 : _GEN_15972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15974 = 7'h3c == _myNewVec_4_T_3[6:0] ? myVec_60 : _GEN_15973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15975 = 7'h3d == _myNewVec_4_T_3[6:0] ? myVec_61 : _GEN_15974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15976 = 7'h3e == _myNewVec_4_T_3[6:0] ? myVec_62 : _GEN_15975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15977 = 7'h3f == _myNewVec_4_T_3[6:0] ? myVec_63 : _GEN_15976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15978 = 7'h40 == _myNewVec_4_T_3[6:0] ? myVec_64 : _GEN_15977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15979 = 7'h41 == _myNewVec_4_T_3[6:0] ? myVec_65 : _GEN_15978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15980 = 7'h42 == _myNewVec_4_T_3[6:0] ? myVec_66 : _GEN_15979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15981 = 7'h43 == _myNewVec_4_T_3[6:0] ? myVec_67 : _GEN_15980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15982 = 7'h44 == _myNewVec_4_T_3[6:0] ? myVec_68 : _GEN_15981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15983 = 7'h45 == _myNewVec_4_T_3[6:0] ? myVec_69 : _GEN_15982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15984 = 7'h46 == _myNewVec_4_T_3[6:0] ? myVec_70 : _GEN_15983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15985 = 7'h47 == _myNewVec_4_T_3[6:0] ? myVec_71 : _GEN_15984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15986 = 7'h48 == _myNewVec_4_T_3[6:0] ? myVec_72 : _GEN_15985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15987 = 7'h49 == _myNewVec_4_T_3[6:0] ? myVec_73 : _GEN_15986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15988 = 7'h4a == _myNewVec_4_T_3[6:0] ? myVec_74 : _GEN_15987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15989 = 7'h4b == _myNewVec_4_T_3[6:0] ? myVec_75 : _GEN_15988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15990 = 7'h4c == _myNewVec_4_T_3[6:0] ? myVec_76 : _GEN_15989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15991 = 7'h4d == _myNewVec_4_T_3[6:0] ? myVec_77 : _GEN_15990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15992 = 7'h4e == _myNewVec_4_T_3[6:0] ? myVec_78 : _GEN_15991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15993 = 7'h4f == _myNewVec_4_T_3[6:0] ? myVec_79 : _GEN_15992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15994 = 7'h50 == _myNewVec_4_T_3[6:0] ? myVec_80 : _GEN_15993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15995 = 7'h51 == _myNewVec_4_T_3[6:0] ? myVec_81 : _GEN_15994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15996 = 7'h52 == _myNewVec_4_T_3[6:0] ? myVec_82 : _GEN_15995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15997 = 7'h53 == _myNewVec_4_T_3[6:0] ? myVec_83 : _GEN_15996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15998 = 7'h54 == _myNewVec_4_T_3[6:0] ? myVec_84 : _GEN_15997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_15999 = 7'h55 == _myNewVec_4_T_3[6:0] ? myVec_85 : _GEN_15998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16000 = 7'h56 == _myNewVec_4_T_3[6:0] ? myVec_86 : _GEN_15999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16001 = 7'h57 == _myNewVec_4_T_3[6:0] ? myVec_87 : _GEN_16000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16002 = 7'h58 == _myNewVec_4_T_3[6:0] ? myVec_88 : _GEN_16001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16003 = 7'h59 == _myNewVec_4_T_3[6:0] ? myVec_89 : _GEN_16002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16004 = 7'h5a == _myNewVec_4_T_3[6:0] ? myVec_90 : _GEN_16003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16005 = 7'h5b == _myNewVec_4_T_3[6:0] ? myVec_91 : _GEN_16004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16006 = 7'h5c == _myNewVec_4_T_3[6:0] ? myVec_92 : _GEN_16005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16007 = 7'h5d == _myNewVec_4_T_3[6:0] ? myVec_93 : _GEN_16006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16008 = 7'h5e == _myNewVec_4_T_3[6:0] ? myVec_94 : _GEN_16007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16009 = 7'h5f == _myNewVec_4_T_3[6:0] ? myVec_95 : _GEN_16008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16010 = 7'h60 == _myNewVec_4_T_3[6:0] ? myVec_96 : _GEN_16009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16011 = 7'h61 == _myNewVec_4_T_3[6:0] ? myVec_97 : _GEN_16010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16012 = 7'h62 == _myNewVec_4_T_3[6:0] ? myVec_98 : _GEN_16011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16013 = 7'h63 == _myNewVec_4_T_3[6:0] ? myVec_99 : _GEN_16012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16014 = 7'h64 == _myNewVec_4_T_3[6:0] ? myVec_100 : _GEN_16013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16015 = 7'h65 == _myNewVec_4_T_3[6:0] ? myVec_101 : _GEN_16014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16016 = 7'h66 == _myNewVec_4_T_3[6:0] ? myVec_102 : _GEN_16015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16017 = 7'h67 == _myNewVec_4_T_3[6:0] ? myVec_103 : _GEN_16016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16018 = 7'h68 == _myNewVec_4_T_3[6:0] ? myVec_104 : _GEN_16017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16019 = 7'h69 == _myNewVec_4_T_3[6:0] ? myVec_105 : _GEN_16018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16020 = 7'h6a == _myNewVec_4_T_3[6:0] ? myVec_106 : _GEN_16019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16021 = 7'h6b == _myNewVec_4_T_3[6:0] ? myVec_107 : _GEN_16020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16022 = 7'h6c == _myNewVec_4_T_3[6:0] ? myVec_108 : _GEN_16021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16023 = 7'h6d == _myNewVec_4_T_3[6:0] ? myVec_109 : _GEN_16022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16024 = 7'h6e == _myNewVec_4_T_3[6:0] ? myVec_110 : _GEN_16023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16025 = 7'h6f == _myNewVec_4_T_3[6:0] ? myVec_111 : _GEN_16024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16026 = 7'h70 == _myNewVec_4_T_3[6:0] ? myVec_112 : _GEN_16025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16027 = 7'h71 == _myNewVec_4_T_3[6:0] ? myVec_113 : _GEN_16026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16028 = 7'h72 == _myNewVec_4_T_3[6:0] ? myVec_114 : _GEN_16027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16029 = 7'h73 == _myNewVec_4_T_3[6:0] ? myVec_115 : _GEN_16028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16030 = 7'h74 == _myNewVec_4_T_3[6:0] ? myVec_116 : _GEN_16029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16031 = 7'h75 == _myNewVec_4_T_3[6:0] ? myVec_117 : _GEN_16030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16032 = 7'h76 == _myNewVec_4_T_3[6:0] ? myVec_118 : _GEN_16031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16033 = 7'h77 == _myNewVec_4_T_3[6:0] ? myVec_119 : _GEN_16032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16034 = 7'h78 == _myNewVec_4_T_3[6:0] ? myVec_120 : _GEN_16033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16035 = 7'h79 == _myNewVec_4_T_3[6:0] ? myVec_121 : _GEN_16034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16036 = 7'h7a == _myNewVec_4_T_3[6:0] ? myVec_122 : _GEN_16035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16037 = 7'h7b == _myNewVec_4_T_3[6:0] ? myVec_123 : _GEN_16036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16038 = 7'h7c == _myNewVec_4_T_3[6:0] ? myVec_124 : _GEN_16037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16039 = 7'h7d == _myNewVec_4_T_3[6:0] ? myVec_125 : _GEN_16038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16040 = 7'h7e == _myNewVec_4_T_3[6:0] ? myVec_126 : _GEN_16039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_4 = 7'h7f == _myNewVec_4_T_3[6:0] ? myVec_127 : _GEN_16040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_3_T_3 = _myNewVec_127_T_1 + 16'h7c; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_16043 = 7'h1 == _myNewVec_3_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16044 = 7'h2 == _myNewVec_3_T_3[6:0] ? myVec_2 : _GEN_16043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16045 = 7'h3 == _myNewVec_3_T_3[6:0] ? myVec_3 : _GEN_16044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16046 = 7'h4 == _myNewVec_3_T_3[6:0] ? myVec_4 : _GEN_16045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16047 = 7'h5 == _myNewVec_3_T_3[6:0] ? myVec_5 : _GEN_16046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16048 = 7'h6 == _myNewVec_3_T_3[6:0] ? myVec_6 : _GEN_16047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16049 = 7'h7 == _myNewVec_3_T_3[6:0] ? myVec_7 : _GEN_16048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16050 = 7'h8 == _myNewVec_3_T_3[6:0] ? myVec_8 : _GEN_16049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16051 = 7'h9 == _myNewVec_3_T_3[6:0] ? myVec_9 : _GEN_16050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16052 = 7'ha == _myNewVec_3_T_3[6:0] ? myVec_10 : _GEN_16051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16053 = 7'hb == _myNewVec_3_T_3[6:0] ? myVec_11 : _GEN_16052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16054 = 7'hc == _myNewVec_3_T_3[6:0] ? myVec_12 : _GEN_16053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16055 = 7'hd == _myNewVec_3_T_3[6:0] ? myVec_13 : _GEN_16054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16056 = 7'he == _myNewVec_3_T_3[6:0] ? myVec_14 : _GEN_16055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16057 = 7'hf == _myNewVec_3_T_3[6:0] ? myVec_15 : _GEN_16056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16058 = 7'h10 == _myNewVec_3_T_3[6:0] ? myVec_16 : _GEN_16057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16059 = 7'h11 == _myNewVec_3_T_3[6:0] ? myVec_17 : _GEN_16058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16060 = 7'h12 == _myNewVec_3_T_3[6:0] ? myVec_18 : _GEN_16059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16061 = 7'h13 == _myNewVec_3_T_3[6:0] ? myVec_19 : _GEN_16060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16062 = 7'h14 == _myNewVec_3_T_3[6:0] ? myVec_20 : _GEN_16061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16063 = 7'h15 == _myNewVec_3_T_3[6:0] ? myVec_21 : _GEN_16062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16064 = 7'h16 == _myNewVec_3_T_3[6:0] ? myVec_22 : _GEN_16063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16065 = 7'h17 == _myNewVec_3_T_3[6:0] ? myVec_23 : _GEN_16064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16066 = 7'h18 == _myNewVec_3_T_3[6:0] ? myVec_24 : _GEN_16065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16067 = 7'h19 == _myNewVec_3_T_3[6:0] ? myVec_25 : _GEN_16066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16068 = 7'h1a == _myNewVec_3_T_3[6:0] ? myVec_26 : _GEN_16067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16069 = 7'h1b == _myNewVec_3_T_3[6:0] ? myVec_27 : _GEN_16068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16070 = 7'h1c == _myNewVec_3_T_3[6:0] ? myVec_28 : _GEN_16069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16071 = 7'h1d == _myNewVec_3_T_3[6:0] ? myVec_29 : _GEN_16070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16072 = 7'h1e == _myNewVec_3_T_3[6:0] ? myVec_30 : _GEN_16071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16073 = 7'h1f == _myNewVec_3_T_3[6:0] ? myVec_31 : _GEN_16072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16074 = 7'h20 == _myNewVec_3_T_3[6:0] ? myVec_32 : _GEN_16073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16075 = 7'h21 == _myNewVec_3_T_3[6:0] ? myVec_33 : _GEN_16074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16076 = 7'h22 == _myNewVec_3_T_3[6:0] ? myVec_34 : _GEN_16075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16077 = 7'h23 == _myNewVec_3_T_3[6:0] ? myVec_35 : _GEN_16076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16078 = 7'h24 == _myNewVec_3_T_3[6:0] ? myVec_36 : _GEN_16077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16079 = 7'h25 == _myNewVec_3_T_3[6:0] ? myVec_37 : _GEN_16078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16080 = 7'h26 == _myNewVec_3_T_3[6:0] ? myVec_38 : _GEN_16079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16081 = 7'h27 == _myNewVec_3_T_3[6:0] ? myVec_39 : _GEN_16080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16082 = 7'h28 == _myNewVec_3_T_3[6:0] ? myVec_40 : _GEN_16081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16083 = 7'h29 == _myNewVec_3_T_3[6:0] ? myVec_41 : _GEN_16082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16084 = 7'h2a == _myNewVec_3_T_3[6:0] ? myVec_42 : _GEN_16083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16085 = 7'h2b == _myNewVec_3_T_3[6:0] ? myVec_43 : _GEN_16084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16086 = 7'h2c == _myNewVec_3_T_3[6:0] ? myVec_44 : _GEN_16085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16087 = 7'h2d == _myNewVec_3_T_3[6:0] ? myVec_45 : _GEN_16086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16088 = 7'h2e == _myNewVec_3_T_3[6:0] ? myVec_46 : _GEN_16087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16089 = 7'h2f == _myNewVec_3_T_3[6:0] ? myVec_47 : _GEN_16088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16090 = 7'h30 == _myNewVec_3_T_3[6:0] ? myVec_48 : _GEN_16089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16091 = 7'h31 == _myNewVec_3_T_3[6:0] ? myVec_49 : _GEN_16090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16092 = 7'h32 == _myNewVec_3_T_3[6:0] ? myVec_50 : _GEN_16091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16093 = 7'h33 == _myNewVec_3_T_3[6:0] ? myVec_51 : _GEN_16092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16094 = 7'h34 == _myNewVec_3_T_3[6:0] ? myVec_52 : _GEN_16093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16095 = 7'h35 == _myNewVec_3_T_3[6:0] ? myVec_53 : _GEN_16094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16096 = 7'h36 == _myNewVec_3_T_3[6:0] ? myVec_54 : _GEN_16095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16097 = 7'h37 == _myNewVec_3_T_3[6:0] ? myVec_55 : _GEN_16096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16098 = 7'h38 == _myNewVec_3_T_3[6:0] ? myVec_56 : _GEN_16097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16099 = 7'h39 == _myNewVec_3_T_3[6:0] ? myVec_57 : _GEN_16098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16100 = 7'h3a == _myNewVec_3_T_3[6:0] ? myVec_58 : _GEN_16099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16101 = 7'h3b == _myNewVec_3_T_3[6:0] ? myVec_59 : _GEN_16100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16102 = 7'h3c == _myNewVec_3_T_3[6:0] ? myVec_60 : _GEN_16101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16103 = 7'h3d == _myNewVec_3_T_3[6:0] ? myVec_61 : _GEN_16102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16104 = 7'h3e == _myNewVec_3_T_3[6:0] ? myVec_62 : _GEN_16103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16105 = 7'h3f == _myNewVec_3_T_3[6:0] ? myVec_63 : _GEN_16104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16106 = 7'h40 == _myNewVec_3_T_3[6:0] ? myVec_64 : _GEN_16105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16107 = 7'h41 == _myNewVec_3_T_3[6:0] ? myVec_65 : _GEN_16106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16108 = 7'h42 == _myNewVec_3_T_3[6:0] ? myVec_66 : _GEN_16107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16109 = 7'h43 == _myNewVec_3_T_3[6:0] ? myVec_67 : _GEN_16108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16110 = 7'h44 == _myNewVec_3_T_3[6:0] ? myVec_68 : _GEN_16109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16111 = 7'h45 == _myNewVec_3_T_3[6:0] ? myVec_69 : _GEN_16110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16112 = 7'h46 == _myNewVec_3_T_3[6:0] ? myVec_70 : _GEN_16111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16113 = 7'h47 == _myNewVec_3_T_3[6:0] ? myVec_71 : _GEN_16112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16114 = 7'h48 == _myNewVec_3_T_3[6:0] ? myVec_72 : _GEN_16113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16115 = 7'h49 == _myNewVec_3_T_3[6:0] ? myVec_73 : _GEN_16114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16116 = 7'h4a == _myNewVec_3_T_3[6:0] ? myVec_74 : _GEN_16115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16117 = 7'h4b == _myNewVec_3_T_3[6:0] ? myVec_75 : _GEN_16116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16118 = 7'h4c == _myNewVec_3_T_3[6:0] ? myVec_76 : _GEN_16117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16119 = 7'h4d == _myNewVec_3_T_3[6:0] ? myVec_77 : _GEN_16118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16120 = 7'h4e == _myNewVec_3_T_3[6:0] ? myVec_78 : _GEN_16119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16121 = 7'h4f == _myNewVec_3_T_3[6:0] ? myVec_79 : _GEN_16120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16122 = 7'h50 == _myNewVec_3_T_3[6:0] ? myVec_80 : _GEN_16121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16123 = 7'h51 == _myNewVec_3_T_3[6:0] ? myVec_81 : _GEN_16122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16124 = 7'h52 == _myNewVec_3_T_3[6:0] ? myVec_82 : _GEN_16123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16125 = 7'h53 == _myNewVec_3_T_3[6:0] ? myVec_83 : _GEN_16124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16126 = 7'h54 == _myNewVec_3_T_3[6:0] ? myVec_84 : _GEN_16125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16127 = 7'h55 == _myNewVec_3_T_3[6:0] ? myVec_85 : _GEN_16126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16128 = 7'h56 == _myNewVec_3_T_3[6:0] ? myVec_86 : _GEN_16127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16129 = 7'h57 == _myNewVec_3_T_3[6:0] ? myVec_87 : _GEN_16128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16130 = 7'h58 == _myNewVec_3_T_3[6:0] ? myVec_88 : _GEN_16129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16131 = 7'h59 == _myNewVec_3_T_3[6:0] ? myVec_89 : _GEN_16130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16132 = 7'h5a == _myNewVec_3_T_3[6:0] ? myVec_90 : _GEN_16131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16133 = 7'h5b == _myNewVec_3_T_3[6:0] ? myVec_91 : _GEN_16132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16134 = 7'h5c == _myNewVec_3_T_3[6:0] ? myVec_92 : _GEN_16133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16135 = 7'h5d == _myNewVec_3_T_3[6:0] ? myVec_93 : _GEN_16134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16136 = 7'h5e == _myNewVec_3_T_3[6:0] ? myVec_94 : _GEN_16135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16137 = 7'h5f == _myNewVec_3_T_3[6:0] ? myVec_95 : _GEN_16136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16138 = 7'h60 == _myNewVec_3_T_3[6:0] ? myVec_96 : _GEN_16137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16139 = 7'h61 == _myNewVec_3_T_3[6:0] ? myVec_97 : _GEN_16138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16140 = 7'h62 == _myNewVec_3_T_3[6:0] ? myVec_98 : _GEN_16139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16141 = 7'h63 == _myNewVec_3_T_3[6:0] ? myVec_99 : _GEN_16140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16142 = 7'h64 == _myNewVec_3_T_3[6:0] ? myVec_100 : _GEN_16141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16143 = 7'h65 == _myNewVec_3_T_3[6:0] ? myVec_101 : _GEN_16142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16144 = 7'h66 == _myNewVec_3_T_3[6:0] ? myVec_102 : _GEN_16143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16145 = 7'h67 == _myNewVec_3_T_3[6:0] ? myVec_103 : _GEN_16144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16146 = 7'h68 == _myNewVec_3_T_3[6:0] ? myVec_104 : _GEN_16145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16147 = 7'h69 == _myNewVec_3_T_3[6:0] ? myVec_105 : _GEN_16146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16148 = 7'h6a == _myNewVec_3_T_3[6:0] ? myVec_106 : _GEN_16147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16149 = 7'h6b == _myNewVec_3_T_3[6:0] ? myVec_107 : _GEN_16148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16150 = 7'h6c == _myNewVec_3_T_3[6:0] ? myVec_108 : _GEN_16149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16151 = 7'h6d == _myNewVec_3_T_3[6:0] ? myVec_109 : _GEN_16150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16152 = 7'h6e == _myNewVec_3_T_3[6:0] ? myVec_110 : _GEN_16151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16153 = 7'h6f == _myNewVec_3_T_3[6:0] ? myVec_111 : _GEN_16152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16154 = 7'h70 == _myNewVec_3_T_3[6:0] ? myVec_112 : _GEN_16153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16155 = 7'h71 == _myNewVec_3_T_3[6:0] ? myVec_113 : _GEN_16154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16156 = 7'h72 == _myNewVec_3_T_3[6:0] ? myVec_114 : _GEN_16155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16157 = 7'h73 == _myNewVec_3_T_3[6:0] ? myVec_115 : _GEN_16156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16158 = 7'h74 == _myNewVec_3_T_3[6:0] ? myVec_116 : _GEN_16157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16159 = 7'h75 == _myNewVec_3_T_3[6:0] ? myVec_117 : _GEN_16158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16160 = 7'h76 == _myNewVec_3_T_3[6:0] ? myVec_118 : _GEN_16159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16161 = 7'h77 == _myNewVec_3_T_3[6:0] ? myVec_119 : _GEN_16160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16162 = 7'h78 == _myNewVec_3_T_3[6:0] ? myVec_120 : _GEN_16161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16163 = 7'h79 == _myNewVec_3_T_3[6:0] ? myVec_121 : _GEN_16162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16164 = 7'h7a == _myNewVec_3_T_3[6:0] ? myVec_122 : _GEN_16163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16165 = 7'h7b == _myNewVec_3_T_3[6:0] ? myVec_123 : _GEN_16164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16166 = 7'h7c == _myNewVec_3_T_3[6:0] ? myVec_124 : _GEN_16165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16167 = 7'h7d == _myNewVec_3_T_3[6:0] ? myVec_125 : _GEN_16166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16168 = 7'h7e == _myNewVec_3_T_3[6:0] ? myVec_126 : _GEN_16167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_3 = 7'h7f == _myNewVec_3_T_3[6:0] ? myVec_127 : _GEN_16168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_2_T_3 = _myNewVec_127_T_1 + 16'h7d; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_16171 = 7'h1 == _myNewVec_2_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16172 = 7'h2 == _myNewVec_2_T_3[6:0] ? myVec_2 : _GEN_16171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16173 = 7'h3 == _myNewVec_2_T_3[6:0] ? myVec_3 : _GEN_16172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16174 = 7'h4 == _myNewVec_2_T_3[6:0] ? myVec_4 : _GEN_16173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16175 = 7'h5 == _myNewVec_2_T_3[6:0] ? myVec_5 : _GEN_16174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16176 = 7'h6 == _myNewVec_2_T_3[6:0] ? myVec_6 : _GEN_16175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16177 = 7'h7 == _myNewVec_2_T_3[6:0] ? myVec_7 : _GEN_16176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16178 = 7'h8 == _myNewVec_2_T_3[6:0] ? myVec_8 : _GEN_16177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16179 = 7'h9 == _myNewVec_2_T_3[6:0] ? myVec_9 : _GEN_16178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16180 = 7'ha == _myNewVec_2_T_3[6:0] ? myVec_10 : _GEN_16179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16181 = 7'hb == _myNewVec_2_T_3[6:0] ? myVec_11 : _GEN_16180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16182 = 7'hc == _myNewVec_2_T_3[6:0] ? myVec_12 : _GEN_16181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16183 = 7'hd == _myNewVec_2_T_3[6:0] ? myVec_13 : _GEN_16182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16184 = 7'he == _myNewVec_2_T_3[6:0] ? myVec_14 : _GEN_16183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16185 = 7'hf == _myNewVec_2_T_3[6:0] ? myVec_15 : _GEN_16184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16186 = 7'h10 == _myNewVec_2_T_3[6:0] ? myVec_16 : _GEN_16185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16187 = 7'h11 == _myNewVec_2_T_3[6:0] ? myVec_17 : _GEN_16186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16188 = 7'h12 == _myNewVec_2_T_3[6:0] ? myVec_18 : _GEN_16187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16189 = 7'h13 == _myNewVec_2_T_3[6:0] ? myVec_19 : _GEN_16188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16190 = 7'h14 == _myNewVec_2_T_3[6:0] ? myVec_20 : _GEN_16189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16191 = 7'h15 == _myNewVec_2_T_3[6:0] ? myVec_21 : _GEN_16190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16192 = 7'h16 == _myNewVec_2_T_3[6:0] ? myVec_22 : _GEN_16191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16193 = 7'h17 == _myNewVec_2_T_3[6:0] ? myVec_23 : _GEN_16192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16194 = 7'h18 == _myNewVec_2_T_3[6:0] ? myVec_24 : _GEN_16193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16195 = 7'h19 == _myNewVec_2_T_3[6:0] ? myVec_25 : _GEN_16194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16196 = 7'h1a == _myNewVec_2_T_3[6:0] ? myVec_26 : _GEN_16195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16197 = 7'h1b == _myNewVec_2_T_3[6:0] ? myVec_27 : _GEN_16196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16198 = 7'h1c == _myNewVec_2_T_3[6:0] ? myVec_28 : _GEN_16197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16199 = 7'h1d == _myNewVec_2_T_3[6:0] ? myVec_29 : _GEN_16198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16200 = 7'h1e == _myNewVec_2_T_3[6:0] ? myVec_30 : _GEN_16199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16201 = 7'h1f == _myNewVec_2_T_3[6:0] ? myVec_31 : _GEN_16200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16202 = 7'h20 == _myNewVec_2_T_3[6:0] ? myVec_32 : _GEN_16201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16203 = 7'h21 == _myNewVec_2_T_3[6:0] ? myVec_33 : _GEN_16202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16204 = 7'h22 == _myNewVec_2_T_3[6:0] ? myVec_34 : _GEN_16203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16205 = 7'h23 == _myNewVec_2_T_3[6:0] ? myVec_35 : _GEN_16204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16206 = 7'h24 == _myNewVec_2_T_3[6:0] ? myVec_36 : _GEN_16205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16207 = 7'h25 == _myNewVec_2_T_3[6:0] ? myVec_37 : _GEN_16206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16208 = 7'h26 == _myNewVec_2_T_3[6:0] ? myVec_38 : _GEN_16207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16209 = 7'h27 == _myNewVec_2_T_3[6:0] ? myVec_39 : _GEN_16208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16210 = 7'h28 == _myNewVec_2_T_3[6:0] ? myVec_40 : _GEN_16209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16211 = 7'h29 == _myNewVec_2_T_3[6:0] ? myVec_41 : _GEN_16210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16212 = 7'h2a == _myNewVec_2_T_3[6:0] ? myVec_42 : _GEN_16211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16213 = 7'h2b == _myNewVec_2_T_3[6:0] ? myVec_43 : _GEN_16212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16214 = 7'h2c == _myNewVec_2_T_3[6:0] ? myVec_44 : _GEN_16213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16215 = 7'h2d == _myNewVec_2_T_3[6:0] ? myVec_45 : _GEN_16214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16216 = 7'h2e == _myNewVec_2_T_3[6:0] ? myVec_46 : _GEN_16215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16217 = 7'h2f == _myNewVec_2_T_3[6:0] ? myVec_47 : _GEN_16216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16218 = 7'h30 == _myNewVec_2_T_3[6:0] ? myVec_48 : _GEN_16217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16219 = 7'h31 == _myNewVec_2_T_3[6:0] ? myVec_49 : _GEN_16218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16220 = 7'h32 == _myNewVec_2_T_3[6:0] ? myVec_50 : _GEN_16219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16221 = 7'h33 == _myNewVec_2_T_3[6:0] ? myVec_51 : _GEN_16220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16222 = 7'h34 == _myNewVec_2_T_3[6:0] ? myVec_52 : _GEN_16221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16223 = 7'h35 == _myNewVec_2_T_3[6:0] ? myVec_53 : _GEN_16222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16224 = 7'h36 == _myNewVec_2_T_3[6:0] ? myVec_54 : _GEN_16223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16225 = 7'h37 == _myNewVec_2_T_3[6:0] ? myVec_55 : _GEN_16224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16226 = 7'h38 == _myNewVec_2_T_3[6:0] ? myVec_56 : _GEN_16225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16227 = 7'h39 == _myNewVec_2_T_3[6:0] ? myVec_57 : _GEN_16226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16228 = 7'h3a == _myNewVec_2_T_3[6:0] ? myVec_58 : _GEN_16227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16229 = 7'h3b == _myNewVec_2_T_3[6:0] ? myVec_59 : _GEN_16228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16230 = 7'h3c == _myNewVec_2_T_3[6:0] ? myVec_60 : _GEN_16229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16231 = 7'h3d == _myNewVec_2_T_3[6:0] ? myVec_61 : _GEN_16230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16232 = 7'h3e == _myNewVec_2_T_3[6:0] ? myVec_62 : _GEN_16231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16233 = 7'h3f == _myNewVec_2_T_3[6:0] ? myVec_63 : _GEN_16232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16234 = 7'h40 == _myNewVec_2_T_3[6:0] ? myVec_64 : _GEN_16233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16235 = 7'h41 == _myNewVec_2_T_3[6:0] ? myVec_65 : _GEN_16234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16236 = 7'h42 == _myNewVec_2_T_3[6:0] ? myVec_66 : _GEN_16235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16237 = 7'h43 == _myNewVec_2_T_3[6:0] ? myVec_67 : _GEN_16236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16238 = 7'h44 == _myNewVec_2_T_3[6:0] ? myVec_68 : _GEN_16237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16239 = 7'h45 == _myNewVec_2_T_3[6:0] ? myVec_69 : _GEN_16238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16240 = 7'h46 == _myNewVec_2_T_3[6:0] ? myVec_70 : _GEN_16239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16241 = 7'h47 == _myNewVec_2_T_3[6:0] ? myVec_71 : _GEN_16240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16242 = 7'h48 == _myNewVec_2_T_3[6:0] ? myVec_72 : _GEN_16241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16243 = 7'h49 == _myNewVec_2_T_3[6:0] ? myVec_73 : _GEN_16242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16244 = 7'h4a == _myNewVec_2_T_3[6:0] ? myVec_74 : _GEN_16243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16245 = 7'h4b == _myNewVec_2_T_3[6:0] ? myVec_75 : _GEN_16244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16246 = 7'h4c == _myNewVec_2_T_3[6:0] ? myVec_76 : _GEN_16245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16247 = 7'h4d == _myNewVec_2_T_3[6:0] ? myVec_77 : _GEN_16246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16248 = 7'h4e == _myNewVec_2_T_3[6:0] ? myVec_78 : _GEN_16247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16249 = 7'h4f == _myNewVec_2_T_3[6:0] ? myVec_79 : _GEN_16248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16250 = 7'h50 == _myNewVec_2_T_3[6:0] ? myVec_80 : _GEN_16249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16251 = 7'h51 == _myNewVec_2_T_3[6:0] ? myVec_81 : _GEN_16250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16252 = 7'h52 == _myNewVec_2_T_3[6:0] ? myVec_82 : _GEN_16251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16253 = 7'h53 == _myNewVec_2_T_3[6:0] ? myVec_83 : _GEN_16252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16254 = 7'h54 == _myNewVec_2_T_3[6:0] ? myVec_84 : _GEN_16253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16255 = 7'h55 == _myNewVec_2_T_3[6:0] ? myVec_85 : _GEN_16254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16256 = 7'h56 == _myNewVec_2_T_3[6:0] ? myVec_86 : _GEN_16255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16257 = 7'h57 == _myNewVec_2_T_3[6:0] ? myVec_87 : _GEN_16256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16258 = 7'h58 == _myNewVec_2_T_3[6:0] ? myVec_88 : _GEN_16257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16259 = 7'h59 == _myNewVec_2_T_3[6:0] ? myVec_89 : _GEN_16258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16260 = 7'h5a == _myNewVec_2_T_3[6:0] ? myVec_90 : _GEN_16259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16261 = 7'h5b == _myNewVec_2_T_3[6:0] ? myVec_91 : _GEN_16260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16262 = 7'h5c == _myNewVec_2_T_3[6:0] ? myVec_92 : _GEN_16261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16263 = 7'h5d == _myNewVec_2_T_3[6:0] ? myVec_93 : _GEN_16262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16264 = 7'h5e == _myNewVec_2_T_3[6:0] ? myVec_94 : _GEN_16263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16265 = 7'h5f == _myNewVec_2_T_3[6:0] ? myVec_95 : _GEN_16264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16266 = 7'h60 == _myNewVec_2_T_3[6:0] ? myVec_96 : _GEN_16265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16267 = 7'h61 == _myNewVec_2_T_3[6:0] ? myVec_97 : _GEN_16266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16268 = 7'h62 == _myNewVec_2_T_3[6:0] ? myVec_98 : _GEN_16267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16269 = 7'h63 == _myNewVec_2_T_3[6:0] ? myVec_99 : _GEN_16268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16270 = 7'h64 == _myNewVec_2_T_3[6:0] ? myVec_100 : _GEN_16269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16271 = 7'h65 == _myNewVec_2_T_3[6:0] ? myVec_101 : _GEN_16270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16272 = 7'h66 == _myNewVec_2_T_3[6:0] ? myVec_102 : _GEN_16271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16273 = 7'h67 == _myNewVec_2_T_3[6:0] ? myVec_103 : _GEN_16272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16274 = 7'h68 == _myNewVec_2_T_3[6:0] ? myVec_104 : _GEN_16273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16275 = 7'h69 == _myNewVec_2_T_3[6:0] ? myVec_105 : _GEN_16274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16276 = 7'h6a == _myNewVec_2_T_3[6:0] ? myVec_106 : _GEN_16275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16277 = 7'h6b == _myNewVec_2_T_3[6:0] ? myVec_107 : _GEN_16276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16278 = 7'h6c == _myNewVec_2_T_3[6:0] ? myVec_108 : _GEN_16277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16279 = 7'h6d == _myNewVec_2_T_3[6:0] ? myVec_109 : _GEN_16278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16280 = 7'h6e == _myNewVec_2_T_3[6:0] ? myVec_110 : _GEN_16279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16281 = 7'h6f == _myNewVec_2_T_3[6:0] ? myVec_111 : _GEN_16280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16282 = 7'h70 == _myNewVec_2_T_3[6:0] ? myVec_112 : _GEN_16281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16283 = 7'h71 == _myNewVec_2_T_3[6:0] ? myVec_113 : _GEN_16282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16284 = 7'h72 == _myNewVec_2_T_3[6:0] ? myVec_114 : _GEN_16283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16285 = 7'h73 == _myNewVec_2_T_3[6:0] ? myVec_115 : _GEN_16284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16286 = 7'h74 == _myNewVec_2_T_3[6:0] ? myVec_116 : _GEN_16285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16287 = 7'h75 == _myNewVec_2_T_3[6:0] ? myVec_117 : _GEN_16286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16288 = 7'h76 == _myNewVec_2_T_3[6:0] ? myVec_118 : _GEN_16287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16289 = 7'h77 == _myNewVec_2_T_3[6:0] ? myVec_119 : _GEN_16288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16290 = 7'h78 == _myNewVec_2_T_3[6:0] ? myVec_120 : _GEN_16289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16291 = 7'h79 == _myNewVec_2_T_3[6:0] ? myVec_121 : _GEN_16290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16292 = 7'h7a == _myNewVec_2_T_3[6:0] ? myVec_122 : _GEN_16291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16293 = 7'h7b == _myNewVec_2_T_3[6:0] ? myVec_123 : _GEN_16292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16294 = 7'h7c == _myNewVec_2_T_3[6:0] ? myVec_124 : _GEN_16293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16295 = 7'h7d == _myNewVec_2_T_3[6:0] ? myVec_125 : _GEN_16294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16296 = 7'h7e == _myNewVec_2_T_3[6:0] ? myVec_126 : _GEN_16295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_2 = 7'h7f == _myNewVec_2_T_3[6:0] ? myVec_127 : _GEN_16296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_1_T_3 = _myNewVec_127_T_1 + 16'h7e; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_16299 = 7'h1 == _myNewVec_1_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16300 = 7'h2 == _myNewVec_1_T_3[6:0] ? myVec_2 : _GEN_16299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16301 = 7'h3 == _myNewVec_1_T_3[6:0] ? myVec_3 : _GEN_16300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16302 = 7'h4 == _myNewVec_1_T_3[6:0] ? myVec_4 : _GEN_16301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16303 = 7'h5 == _myNewVec_1_T_3[6:0] ? myVec_5 : _GEN_16302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16304 = 7'h6 == _myNewVec_1_T_3[6:0] ? myVec_6 : _GEN_16303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16305 = 7'h7 == _myNewVec_1_T_3[6:0] ? myVec_7 : _GEN_16304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16306 = 7'h8 == _myNewVec_1_T_3[6:0] ? myVec_8 : _GEN_16305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16307 = 7'h9 == _myNewVec_1_T_3[6:0] ? myVec_9 : _GEN_16306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16308 = 7'ha == _myNewVec_1_T_3[6:0] ? myVec_10 : _GEN_16307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16309 = 7'hb == _myNewVec_1_T_3[6:0] ? myVec_11 : _GEN_16308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16310 = 7'hc == _myNewVec_1_T_3[6:0] ? myVec_12 : _GEN_16309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16311 = 7'hd == _myNewVec_1_T_3[6:0] ? myVec_13 : _GEN_16310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16312 = 7'he == _myNewVec_1_T_3[6:0] ? myVec_14 : _GEN_16311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16313 = 7'hf == _myNewVec_1_T_3[6:0] ? myVec_15 : _GEN_16312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16314 = 7'h10 == _myNewVec_1_T_3[6:0] ? myVec_16 : _GEN_16313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16315 = 7'h11 == _myNewVec_1_T_3[6:0] ? myVec_17 : _GEN_16314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16316 = 7'h12 == _myNewVec_1_T_3[6:0] ? myVec_18 : _GEN_16315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16317 = 7'h13 == _myNewVec_1_T_3[6:0] ? myVec_19 : _GEN_16316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16318 = 7'h14 == _myNewVec_1_T_3[6:0] ? myVec_20 : _GEN_16317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16319 = 7'h15 == _myNewVec_1_T_3[6:0] ? myVec_21 : _GEN_16318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16320 = 7'h16 == _myNewVec_1_T_3[6:0] ? myVec_22 : _GEN_16319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16321 = 7'h17 == _myNewVec_1_T_3[6:0] ? myVec_23 : _GEN_16320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16322 = 7'h18 == _myNewVec_1_T_3[6:0] ? myVec_24 : _GEN_16321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16323 = 7'h19 == _myNewVec_1_T_3[6:0] ? myVec_25 : _GEN_16322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16324 = 7'h1a == _myNewVec_1_T_3[6:0] ? myVec_26 : _GEN_16323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16325 = 7'h1b == _myNewVec_1_T_3[6:0] ? myVec_27 : _GEN_16324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16326 = 7'h1c == _myNewVec_1_T_3[6:0] ? myVec_28 : _GEN_16325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16327 = 7'h1d == _myNewVec_1_T_3[6:0] ? myVec_29 : _GEN_16326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16328 = 7'h1e == _myNewVec_1_T_3[6:0] ? myVec_30 : _GEN_16327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16329 = 7'h1f == _myNewVec_1_T_3[6:0] ? myVec_31 : _GEN_16328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16330 = 7'h20 == _myNewVec_1_T_3[6:0] ? myVec_32 : _GEN_16329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16331 = 7'h21 == _myNewVec_1_T_3[6:0] ? myVec_33 : _GEN_16330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16332 = 7'h22 == _myNewVec_1_T_3[6:0] ? myVec_34 : _GEN_16331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16333 = 7'h23 == _myNewVec_1_T_3[6:0] ? myVec_35 : _GEN_16332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16334 = 7'h24 == _myNewVec_1_T_3[6:0] ? myVec_36 : _GEN_16333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16335 = 7'h25 == _myNewVec_1_T_3[6:0] ? myVec_37 : _GEN_16334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16336 = 7'h26 == _myNewVec_1_T_3[6:0] ? myVec_38 : _GEN_16335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16337 = 7'h27 == _myNewVec_1_T_3[6:0] ? myVec_39 : _GEN_16336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16338 = 7'h28 == _myNewVec_1_T_3[6:0] ? myVec_40 : _GEN_16337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16339 = 7'h29 == _myNewVec_1_T_3[6:0] ? myVec_41 : _GEN_16338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16340 = 7'h2a == _myNewVec_1_T_3[6:0] ? myVec_42 : _GEN_16339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16341 = 7'h2b == _myNewVec_1_T_3[6:0] ? myVec_43 : _GEN_16340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16342 = 7'h2c == _myNewVec_1_T_3[6:0] ? myVec_44 : _GEN_16341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16343 = 7'h2d == _myNewVec_1_T_3[6:0] ? myVec_45 : _GEN_16342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16344 = 7'h2e == _myNewVec_1_T_3[6:0] ? myVec_46 : _GEN_16343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16345 = 7'h2f == _myNewVec_1_T_3[6:0] ? myVec_47 : _GEN_16344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16346 = 7'h30 == _myNewVec_1_T_3[6:0] ? myVec_48 : _GEN_16345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16347 = 7'h31 == _myNewVec_1_T_3[6:0] ? myVec_49 : _GEN_16346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16348 = 7'h32 == _myNewVec_1_T_3[6:0] ? myVec_50 : _GEN_16347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16349 = 7'h33 == _myNewVec_1_T_3[6:0] ? myVec_51 : _GEN_16348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16350 = 7'h34 == _myNewVec_1_T_3[6:0] ? myVec_52 : _GEN_16349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16351 = 7'h35 == _myNewVec_1_T_3[6:0] ? myVec_53 : _GEN_16350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16352 = 7'h36 == _myNewVec_1_T_3[6:0] ? myVec_54 : _GEN_16351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16353 = 7'h37 == _myNewVec_1_T_3[6:0] ? myVec_55 : _GEN_16352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16354 = 7'h38 == _myNewVec_1_T_3[6:0] ? myVec_56 : _GEN_16353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16355 = 7'h39 == _myNewVec_1_T_3[6:0] ? myVec_57 : _GEN_16354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16356 = 7'h3a == _myNewVec_1_T_3[6:0] ? myVec_58 : _GEN_16355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16357 = 7'h3b == _myNewVec_1_T_3[6:0] ? myVec_59 : _GEN_16356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16358 = 7'h3c == _myNewVec_1_T_3[6:0] ? myVec_60 : _GEN_16357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16359 = 7'h3d == _myNewVec_1_T_3[6:0] ? myVec_61 : _GEN_16358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16360 = 7'h3e == _myNewVec_1_T_3[6:0] ? myVec_62 : _GEN_16359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16361 = 7'h3f == _myNewVec_1_T_3[6:0] ? myVec_63 : _GEN_16360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16362 = 7'h40 == _myNewVec_1_T_3[6:0] ? myVec_64 : _GEN_16361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16363 = 7'h41 == _myNewVec_1_T_3[6:0] ? myVec_65 : _GEN_16362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16364 = 7'h42 == _myNewVec_1_T_3[6:0] ? myVec_66 : _GEN_16363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16365 = 7'h43 == _myNewVec_1_T_3[6:0] ? myVec_67 : _GEN_16364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16366 = 7'h44 == _myNewVec_1_T_3[6:0] ? myVec_68 : _GEN_16365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16367 = 7'h45 == _myNewVec_1_T_3[6:0] ? myVec_69 : _GEN_16366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16368 = 7'h46 == _myNewVec_1_T_3[6:0] ? myVec_70 : _GEN_16367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16369 = 7'h47 == _myNewVec_1_T_3[6:0] ? myVec_71 : _GEN_16368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16370 = 7'h48 == _myNewVec_1_T_3[6:0] ? myVec_72 : _GEN_16369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16371 = 7'h49 == _myNewVec_1_T_3[6:0] ? myVec_73 : _GEN_16370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16372 = 7'h4a == _myNewVec_1_T_3[6:0] ? myVec_74 : _GEN_16371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16373 = 7'h4b == _myNewVec_1_T_3[6:0] ? myVec_75 : _GEN_16372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16374 = 7'h4c == _myNewVec_1_T_3[6:0] ? myVec_76 : _GEN_16373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16375 = 7'h4d == _myNewVec_1_T_3[6:0] ? myVec_77 : _GEN_16374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16376 = 7'h4e == _myNewVec_1_T_3[6:0] ? myVec_78 : _GEN_16375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16377 = 7'h4f == _myNewVec_1_T_3[6:0] ? myVec_79 : _GEN_16376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16378 = 7'h50 == _myNewVec_1_T_3[6:0] ? myVec_80 : _GEN_16377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16379 = 7'h51 == _myNewVec_1_T_3[6:0] ? myVec_81 : _GEN_16378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16380 = 7'h52 == _myNewVec_1_T_3[6:0] ? myVec_82 : _GEN_16379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16381 = 7'h53 == _myNewVec_1_T_3[6:0] ? myVec_83 : _GEN_16380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16382 = 7'h54 == _myNewVec_1_T_3[6:0] ? myVec_84 : _GEN_16381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16383 = 7'h55 == _myNewVec_1_T_3[6:0] ? myVec_85 : _GEN_16382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16384 = 7'h56 == _myNewVec_1_T_3[6:0] ? myVec_86 : _GEN_16383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16385 = 7'h57 == _myNewVec_1_T_3[6:0] ? myVec_87 : _GEN_16384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16386 = 7'h58 == _myNewVec_1_T_3[6:0] ? myVec_88 : _GEN_16385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16387 = 7'h59 == _myNewVec_1_T_3[6:0] ? myVec_89 : _GEN_16386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16388 = 7'h5a == _myNewVec_1_T_3[6:0] ? myVec_90 : _GEN_16387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16389 = 7'h5b == _myNewVec_1_T_3[6:0] ? myVec_91 : _GEN_16388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16390 = 7'h5c == _myNewVec_1_T_3[6:0] ? myVec_92 : _GEN_16389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16391 = 7'h5d == _myNewVec_1_T_3[6:0] ? myVec_93 : _GEN_16390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16392 = 7'h5e == _myNewVec_1_T_3[6:0] ? myVec_94 : _GEN_16391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16393 = 7'h5f == _myNewVec_1_T_3[6:0] ? myVec_95 : _GEN_16392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16394 = 7'h60 == _myNewVec_1_T_3[6:0] ? myVec_96 : _GEN_16393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16395 = 7'h61 == _myNewVec_1_T_3[6:0] ? myVec_97 : _GEN_16394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16396 = 7'h62 == _myNewVec_1_T_3[6:0] ? myVec_98 : _GEN_16395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16397 = 7'h63 == _myNewVec_1_T_3[6:0] ? myVec_99 : _GEN_16396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16398 = 7'h64 == _myNewVec_1_T_3[6:0] ? myVec_100 : _GEN_16397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16399 = 7'h65 == _myNewVec_1_T_3[6:0] ? myVec_101 : _GEN_16398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16400 = 7'h66 == _myNewVec_1_T_3[6:0] ? myVec_102 : _GEN_16399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16401 = 7'h67 == _myNewVec_1_T_3[6:0] ? myVec_103 : _GEN_16400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16402 = 7'h68 == _myNewVec_1_T_3[6:0] ? myVec_104 : _GEN_16401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16403 = 7'h69 == _myNewVec_1_T_3[6:0] ? myVec_105 : _GEN_16402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16404 = 7'h6a == _myNewVec_1_T_3[6:0] ? myVec_106 : _GEN_16403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16405 = 7'h6b == _myNewVec_1_T_3[6:0] ? myVec_107 : _GEN_16404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16406 = 7'h6c == _myNewVec_1_T_3[6:0] ? myVec_108 : _GEN_16405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16407 = 7'h6d == _myNewVec_1_T_3[6:0] ? myVec_109 : _GEN_16406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16408 = 7'h6e == _myNewVec_1_T_3[6:0] ? myVec_110 : _GEN_16407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16409 = 7'h6f == _myNewVec_1_T_3[6:0] ? myVec_111 : _GEN_16408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16410 = 7'h70 == _myNewVec_1_T_3[6:0] ? myVec_112 : _GEN_16409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16411 = 7'h71 == _myNewVec_1_T_3[6:0] ? myVec_113 : _GEN_16410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16412 = 7'h72 == _myNewVec_1_T_3[6:0] ? myVec_114 : _GEN_16411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16413 = 7'h73 == _myNewVec_1_T_3[6:0] ? myVec_115 : _GEN_16412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16414 = 7'h74 == _myNewVec_1_T_3[6:0] ? myVec_116 : _GEN_16413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16415 = 7'h75 == _myNewVec_1_T_3[6:0] ? myVec_117 : _GEN_16414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16416 = 7'h76 == _myNewVec_1_T_3[6:0] ? myVec_118 : _GEN_16415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16417 = 7'h77 == _myNewVec_1_T_3[6:0] ? myVec_119 : _GEN_16416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16418 = 7'h78 == _myNewVec_1_T_3[6:0] ? myVec_120 : _GEN_16417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16419 = 7'h79 == _myNewVec_1_T_3[6:0] ? myVec_121 : _GEN_16418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16420 = 7'h7a == _myNewVec_1_T_3[6:0] ? myVec_122 : _GEN_16419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16421 = 7'h7b == _myNewVec_1_T_3[6:0] ? myVec_123 : _GEN_16420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16422 = 7'h7c == _myNewVec_1_T_3[6:0] ? myVec_124 : _GEN_16421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16423 = 7'h7d == _myNewVec_1_T_3[6:0] ? myVec_125 : _GEN_16422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16424 = 7'h7e == _myNewVec_1_T_3[6:0] ? myVec_126 : _GEN_16423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_1 = 7'h7f == _myNewVec_1_T_3[6:0] ? myVec_127 : _GEN_16424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_0_T_3 = _myNewVec_127_T_1 + 16'h7f; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_16427 = 7'h1 == _myNewVec_0_T_3[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16428 = 7'h2 == _myNewVec_0_T_3[6:0] ? myVec_2 : _GEN_16427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16429 = 7'h3 == _myNewVec_0_T_3[6:0] ? myVec_3 : _GEN_16428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16430 = 7'h4 == _myNewVec_0_T_3[6:0] ? myVec_4 : _GEN_16429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16431 = 7'h5 == _myNewVec_0_T_3[6:0] ? myVec_5 : _GEN_16430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16432 = 7'h6 == _myNewVec_0_T_3[6:0] ? myVec_6 : _GEN_16431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16433 = 7'h7 == _myNewVec_0_T_3[6:0] ? myVec_7 : _GEN_16432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16434 = 7'h8 == _myNewVec_0_T_3[6:0] ? myVec_8 : _GEN_16433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16435 = 7'h9 == _myNewVec_0_T_3[6:0] ? myVec_9 : _GEN_16434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16436 = 7'ha == _myNewVec_0_T_3[6:0] ? myVec_10 : _GEN_16435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16437 = 7'hb == _myNewVec_0_T_3[6:0] ? myVec_11 : _GEN_16436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16438 = 7'hc == _myNewVec_0_T_3[6:0] ? myVec_12 : _GEN_16437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16439 = 7'hd == _myNewVec_0_T_3[6:0] ? myVec_13 : _GEN_16438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16440 = 7'he == _myNewVec_0_T_3[6:0] ? myVec_14 : _GEN_16439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16441 = 7'hf == _myNewVec_0_T_3[6:0] ? myVec_15 : _GEN_16440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16442 = 7'h10 == _myNewVec_0_T_3[6:0] ? myVec_16 : _GEN_16441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16443 = 7'h11 == _myNewVec_0_T_3[6:0] ? myVec_17 : _GEN_16442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16444 = 7'h12 == _myNewVec_0_T_3[6:0] ? myVec_18 : _GEN_16443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16445 = 7'h13 == _myNewVec_0_T_3[6:0] ? myVec_19 : _GEN_16444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16446 = 7'h14 == _myNewVec_0_T_3[6:0] ? myVec_20 : _GEN_16445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16447 = 7'h15 == _myNewVec_0_T_3[6:0] ? myVec_21 : _GEN_16446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16448 = 7'h16 == _myNewVec_0_T_3[6:0] ? myVec_22 : _GEN_16447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16449 = 7'h17 == _myNewVec_0_T_3[6:0] ? myVec_23 : _GEN_16448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16450 = 7'h18 == _myNewVec_0_T_3[6:0] ? myVec_24 : _GEN_16449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16451 = 7'h19 == _myNewVec_0_T_3[6:0] ? myVec_25 : _GEN_16450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16452 = 7'h1a == _myNewVec_0_T_3[6:0] ? myVec_26 : _GEN_16451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16453 = 7'h1b == _myNewVec_0_T_3[6:0] ? myVec_27 : _GEN_16452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16454 = 7'h1c == _myNewVec_0_T_3[6:0] ? myVec_28 : _GEN_16453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16455 = 7'h1d == _myNewVec_0_T_3[6:0] ? myVec_29 : _GEN_16454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16456 = 7'h1e == _myNewVec_0_T_3[6:0] ? myVec_30 : _GEN_16455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16457 = 7'h1f == _myNewVec_0_T_3[6:0] ? myVec_31 : _GEN_16456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16458 = 7'h20 == _myNewVec_0_T_3[6:0] ? myVec_32 : _GEN_16457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16459 = 7'h21 == _myNewVec_0_T_3[6:0] ? myVec_33 : _GEN_16458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16460 = 7'h22 == _myNewVec_0_T_3[6:0] ? myVec_34 : _GEN_16459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16461 = 7'h23 == _myNewVec_0_T_3[6:0] ? myVec_35 : _GEN_16460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16462 = 7'h24 == _myNewVec_0_T_3[6:0] ? myVec_36 : _GEN_16461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16463 = 7'h25 == _myNewVec_0_T_3[6:0] ? myVec_37 : _GEN_16462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16464 = 7'h26 == _myNewVec_0_T_3[6:0] ? myVec_38 : _GEN_16463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16465 = 7'h27 == _myNewVec_0_T_3[6:0] ? myVec_39 : _GEN_16464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16466 = 7'h28 == _myNewVec_0_T_3[6:0] ? myVec_40 : _GEN_16465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16467 = 7'h29 == _myNewVec_0_T_3[6:0] ? myVec_41 : _GEN_16466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16468 = 7'h2a == _myNewVec_0_T_3[6:0] ? myVec_42 : _GEN_16467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16469 = 7'h2b == _myNewVec_0_T_3[6:0] ? myVec_43 : _GEN_16468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16470 = 7'h2c == _myNewVec_0_T_3[6:0] ? myVec_44 : _GEN_16469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16471 = 7'h2d == _myNewVec_0_T_3[6:0] ? myVec_45 : _GEN_16470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16472 = 7'h2e == _myNewVec_0_T_3[6:0] ? myVec_46 : _GEN_16471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16473 = 7'h2f == _myNewVec_0_T_3[6:0] ? myVec_47 : _GEN_16472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16474 = 7'h30 == _myNewVec_0_T_3[6:0] ? myVec_48 : _GEN_16473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16475 = 7'h31 == _myNewVec_0_T_3[6:0] ? myVec_49 : _GEN_16474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16476 = 7'h32 == _myNewVec_0_T_3[6:0] ? myVec_50 : _GEN_16475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16477 = 7'h33 == _myNewVec_0_T_3[6:0] ? myVec_51 : _GEN_16476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16478 = 7'h34 == _myNewVec_0_T_3[6:0] ? myVec_52 : _GEN_16477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16479 = 7'h35 == _myNewVec_0_T_3[6:0] ? myVec_53 : _GEN_16478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16480 = 7'h36 == _myNewVec_0_T_3[6:0] ? myVec_54 : _GEN_16479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16481 = 7'h37 == _myNewVec_0_T_3[6:0] ? myVec_55 : _GEN_16480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16482 = 7'h38 == _myNewVec_0_T_3[6:0] ? myVec_56 : _GEN_16481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16483 = 7'h39 == _myNewVec_0_T_3[6:0] ? myVec_57 : _GEN_16482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16484 = 7'h3a == _myNewVec_0_T_3[6:0] ? myVec_58 : _GEN_16483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16485 = 7'h3b == _myNewVec_0_T_3[6:0] ? myVec_59 : _GEN_16484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16486 = 7'h3c == _myNewVec_0_T_3[6:0] ? myVec_60 : _GEN_16485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16487 = 7'h3d == _myNewVec_0_T_3[6:0] ? myVec_61 : _GEN_16486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16488 = 7'h3e == _myNewVec_0_T_3[6:0] ? myVec_62 : _GEN_16487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16489 = 7'h3f == _myNewVec_0_T_3[6:0] ? myVec_63 : _GEN_16488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16490 = 7'h40 == _myNewVec_0_T_3[6:0] ? myVec_64 : _GEN_16489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16491 = 7'h41 == _myNewVec_0_T_3[6:0] ? myVec_65 : _GEN_16490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16492 = 7'h42 == _myNewVec_0_T_3[6:0] ? myVec_66 : _GEN_16491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16493 = 7'h43 == _myNewVec_0_T_3[6:0] ? myVec_67 : _GEN_16492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16494 = 7'h44 == _myNewVec_0_T_3[6:0] ? myVec_68 : _GEN_16493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16495 = 7'h45 == _myNewVec_0_T_3[6:0] ? myVec_69 : _GEN_16494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16496 = 7'h46 == _myNewVec_0_T_3[6:0] ? myVec_70 : _GEN_16495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16497 = 7'h47 == _myNewVec_0_T_3[6:0] ? myVec_71 : _GEN_16496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16498 = 7'h48 == _myNewVec_0_T_3[6:0] ? myVec_72 : _GEN_16497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16499 = 7'h49 == _myNewVec_0_T_3[6:0] ? myVec_73 : _GEN_16498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16500 = 7'h4a == _myNewVec_0_T_3[6:0] ? myVec_74 : _GEN_16499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16501 = 7'h4b == _myNewVec_0_T_3[6:0] ? myVec_75 : _GEN_16500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16502 = 7'h4c == _myNewVec_0_T_3[6:0] ? myVec_76 : _GEN_16501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16503 = 7'h4d == _myNewVec_0_T_3[6:0] ? myVec_77 : _GEN_16502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16504 = 7'h4e == _myNewVec_0_T_3[6:0] ? myVec_78 : _GEN_16503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16505 = 7'h4f == _myNewVec_0_T_3[6:0] ? myVec_79 : _GEN_16504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16506 = 7'h50 == _myNewVec_0_T_3[6:0] ? myVec_80 : _GEN_16505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16507 = 7'h51 == _myNewVec_0_T_3[6:0] ? myVec_81 : _GEN_16506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16508 = 7'h52 == _myNewVec_0_T_3[6:0] ? myVec_82 : _GEN_16507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16509 = 7'h53 == _myNewVec_0_T_3[6:0] ? myVec_83 : _GEN_16508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16510 = 7'h54 == _myNewVec_0_T_3[6:0] ? myVec_84 : _GEN_16509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16511 = 7'h55 == _myNewVec_0_T_3[6:0] ? myVec_85 : _GEN_16510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16512 = 7'h56 == _myNewVec_0_T_3[6:0] ? myVec_86 : _GEN_16511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16513 = 7'h57 == _myNewVec_0_T_3[6:0] ? myVec_87 : _GEN_16512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16514 = 7'h58 == _myNewVec_0_T_3[6:0] ? myVec_88 : _GEN_16513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16515 = 7'h59 == _myNewVec_0_T_3[6:0] ? myVec_89 : _GEN_16514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16516 = 7'h5a == _myNewVec_0_T_3[6:0] ? myVec_90 : _GEN_16515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16517 = 7'h5b == _myNewVec_0_T_3[6:0] ? myVec_91 : _GEN_16516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16518 = 7'h5c == _myNewVec_0_T_3[6:0] ? myVec_92 : _GEN_16517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16519 = 7'h5d == _myNewVec_0_T_3[6:0] ? myVec_93 : _GEN_16518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16520 = 7'h5e == _myNewVec_0_T_3[6:0] ? myVec_94 : _GEN_16519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16521 = 7'h5f == _myNewVec_0_T_3[6:0] ? myVec_95 : _GEN_16520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16522 = 7'h60 == _myNewVec_0_T_3[6:0] ? myVec_96 : _GEN_16521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16523 = 7'h61 == _myNewVec_0_T_3[6:0] ? myVec_97 : _GEN_16522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16524 = 7'h62 == _myNewVec_0_T_3[6:0] ? myVec_98 : _GEN_16523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16525 = 7'h63 == _myNewVec_0_T_3[6:0] ? myVec_99 : _GEN_16524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16526 = 7'h64 == _myNewVec_0_T_3[6:0] ? myVec_100 : _GEN_16525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16527 = 7'h65 == _myNewVec_0_T_3[6:0] ? myVec_101 : _GEN_16526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16528 = 7'h66 == _myNewVec_0_T_3[6:0] ? myVec_102 : _GEN_16527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16529 = 7'h67 == _myNewVec_0_T_3[6:0] ? myVec_103 : _GEN_16528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16530 = 7'h68 == _myNewVec_0_T_3[6:0] ? myVec_104 : _GEN_16529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16531 = 7'h69 == _myNewVec_0_T_3[6:0] ? myVec_105 : _GEN_16530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16532 = 7'h6a == _myNewVec_0_T_3[6:0] ? myVec_106 : _GEN_16531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16533 = 7'h6b == _myNewVec_0_T_3[6:0] ? myVec_107 : _GEN_16532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16534 = 7'h6c == _myNewVec_0_T_3[6:0] ? myVec_108 : _GEN_16533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16535 = 7'h6d == _myNewVec_0_T_3[6:0] ? myVec_109 : _GEN_16534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16536 = 7'h6e == _myNewVec_0_T_3[6:0] ? myVec_110 : _GEN_16535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16537 = 7'h6f == _myNewVec_0_T_3[6:0] ? myVec_111 : _GEN_16536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16538 = 7'h70 == _myNewVec_0_T_3[6:0] ? myVec_112 : _GEN_16537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16539 = 7'h71 == _myNewVec_0_T_3[6:0] ? myVec_113 : _GEN_16538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16540 = 7'h72 == _myNewVec_0_T_3[6:0] ? myVec_114 : _GEN_16539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16541 = 7'h73 == _myNewVec_0_T_3[6:0] ? myVec_115 : _GEN_16540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16542 = 7'h74 == _myNewVec_0_T_3[6:0] ? myVec_116 : _GEN_16541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16543 = 7'h75 == _myNewVec_0_T_3[6:0] ? myVec_117 : _GEN_16542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16544 = 7'h76 == _myNewVec_0_T_3[6:0] ? myVec_118 : _GEN_16543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16545 = 7'h77 == _myNewVec_0_T_3[6:0] ? myVec_119 : _GEN_16544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16546 = 7'h78 == _myNewVec_0_T_3[6:0] ? myVec_120 : _GEN_16545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16547 = 7'h79 == _myNewVec_0_T_3[6:0] ? myVec_121 : _GEN_16546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16548 = 7'h7a == _myNewVec_0_T_3[6:0] ? myVec_122 : _GEN_16547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16549 = 7'h7b == _myNewVec_0_T_3[6:0] ? myVec_123 : _GEN_16548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16550 = 7'h7c == _myNewVec_0_T_3[6:0] ? myVec_124 : _GEN_16549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16551 = 7'h7d == _myNewVec_0_T_3[6:0] ? myVec_125 : _GEN_16550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_16552 = 7'h7e == _myNewVec_0_T_3[6:0] ? myVec_126 : _GEN_16551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_0 = 7'h7f == _myNewVec_0_T_3[6:0] ? myVec_127 : _GEN_16552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [255:0] myNewWire_lo_lo_lo_lo = {myNewVec_7,myNewVec_6,myNewVec_5,myNewVec_4,myNewVec_3,myNewVec_2,myNewVec_1,
    myNewVec_0}; // @[hh_datapath_chisel.scala 238:27]
  wire [511:0] myNewWire_lo_lo_lo = {myNewVec_15,myNewVec_14,myNewVec_13,myNewVec_12,myNewVec_11,myNewVec_10,myNewVec_9,
    myNewVec_8,myNewWire_lo_lo_lo_lo}; // @[hh_datapath_chisel.scala 238:27]
  wire [1023:0] myNewWire_lo_lo = {myNewVec_31,myNewVec_30,myNewVec_29,myNewVec_28,myNewVec_27,myNewVec_26,myNewVec_25,
    myNewVec_24,myNewWire_lo_lo_hi_lo,myNewWire_lo_lo_lo}; // @[hh_datapath_chisel.scala 238:27]
  wire [4127:0] _vk_update_T = {vk1,myNewWire_hi_hi,myNewWire_hi_lo,myNewWire_lo_hi,myNewWire_lo_lo}; // @[Cat.scala 31:58]
  wire [21:0] _vk_update_T_3 = _myNewVec_127_T_1 * 6'h20; // @[hh_datapath_chisel.scala 242:57]
  wire [4127:0] _vk_update_T_4 = _vk_update_T >> _vk_update_T_3; // @[hh_datapath_chisel.scala 242:39]
  wire [4127:0] _GEN_16554 = io_vk1_vld ? _vk_update_T_4 : 4128'h0; // @[hh_datapath_chisel.scala 241:27 242:17 245:17]
  wire [4127:0] _GEN_16555 = io_rst ? 4128'h0 : _GEN_16554; // @[hh_datapath_chisel.scala 239:17 240:17]
  wire [4095:0] vk_update = _GEN_16555[4095:0]; // @[hh_datapath_chisel.scala 81:25]
  wire [4095:0] vk = io_vk1_vld ? vk_update : vk_reg; // @[hh_datapath_chisel.scala 155:21 156:10 158:10]
  wire [4095:0] _GEN_21 = io_d4_rdy ? io_hh_din : ddot_din_a_reg; // @[hh_datapath_chisel.scala 139:26 140:18 142:18]
  wire [4095:0] _GEN_22 = io_d3_rdy ? vk : _GEN_21; // @[hh_datapath_chisel.scala 137:26 138:18]
  wire [4095:0] ddot_din_a = io_d1_rdy ? io_hh_din : _GEN_22; // @[hh_datapath_chisel.scala 135:20 136:18]
  wire [4095:0] _GEN_24 = io_d4_rdy ? vk : ddot_din_b_reg; // @[hh_datapath_chisel.scala 149:26 150:18 152:18]
  wire [4095:0] _GEN_25 = io_d3_rdy ? vk : _GEN_24; // @[hh_datapath_chisel.scala 147:26 148:18]
  wire [4095:0] ddot_din_b = io_d1_rdy ? io_hh_din : _GEN_25; // @[hh_datapath_chisel.scala 145:20 146:18]
  wire [31:0] ddot_dout = FP_DDOT_dp_io_out_s; // @[hh_datapath_chisel.scala 254:15 75:25]
  wire [31:0] _GEN_41 = 7'h1 == io_hh_cnt[6:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_42 = 7'h2 == io_hh_cnt[6:0] ? myVec_2 : _GEN_41; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_43 = 7'h3 == io_hh_cnt[6:0] ? myVec_3 : _GEN_42; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_44 = 7'h4 == io_hh_cnt[6:0] ? myVec_4 : _GEN_43; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_45 = 7'h5 == io_hh_cnt[6:0] ? myVec_5 : _GEN_44; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_46 = 7'h6 == io_hh_cnt[6:0] ? myVec_6 : _GEN_45; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_47 = 7'h7 == io_hh_cnt[6:0] ? myVec_7 : _GEN_46; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_48 = 7'h8 == io_hh_cnt[6:0] ? myVec_8 : _GEN_47; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_49 = 7'h9 == io_hh_cnt[6:0] ? myVec_9 : _GEN_48; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_50 = 7'ha == io_hh_cnt[6:0] ? myVec_10 : _GEN_49; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_51 = 7'hb == io_hh_cnt[6:0] ? myVec_11 : _GEN_50; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_52 = 7'hc == io_hh_cnt[6:0] ? myVec_12 : _GEN_51; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_53 = 7'hd == io_hh_cnt[6:0] ? myVec_13 : _GEN_52; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_54 = 7'he == io_hh_cnt[6:0] ? myVec_14 : _GEN_53; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_55 = 7'hf == io_hh_cnt[6:0] ? myVec_15 : _GEN_54; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_56 = 7'h10 == io_hh_cnt[6:0] ? myVec_16 : _GEN_55; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_57 = 7'h11 == io_hh_cnt[6:0] ? myVec_17 : _GEN_56; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_58 = 7'h12 == io_hh_cnt[6:0] ? myVec_18 : _GEN_57; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_59 = 7'h13 == io_hh_cnt[6:0] ? myVec_19 : _GEN_58; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_60 = 7'h14 == io_hh_cnt[6:0] ? myVec_20 : _GEN_59; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_61 = 7'h15 == io_hh_cnt[6:0] ? myVec_21 : _GEN_60; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_62 = 7'h16 == io_hh_cnt[6:0] ? myVec_22 : _GEN_61; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_63 = 7'h17 == io_hh_cnt[6:0] ? myVec_23 : _GEN_62; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_64 = 7'h18 == io_hh_cnt[6:0] ? myVec_24 : _GEN_63; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_65 = 7'h19 == io_hh_cnt[6:0] ? myVec_25 : _GEN_64; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_66 = 7'h1a == io_hh_cnt[6:0] ? myVec_26 : _GEN_65; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_67 = 7'h1b == io_hh_cnt[6:0] ? myVec_27 : _GEN_66; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_68 = 7'h1c == io_hh_cnt[6:0] ? myVec_28 : _GEN_67; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_69 = 7'h1d == io_hh_cnt[6:0] ? myVec_29 : _GEN_68; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_70 = 7'h1e == io_hh_cnt[6:0] ? myVec_30 : _GEN_69; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_71 = 7'h1f == io_hh_cnt[6:0] ? myVec_31 : _GEN_70; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_72 = 7'h20 == io_hh_cnt[6:0] ? myVec_32 : _GEN_71; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_73 = 7'h21 == io_hh_cnt[6:0] ? myVec_33 : _GEN_72; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_74 = 7'h22 == io_hh_cnt[6:0] ? myVec_34 : _GEN_73; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_75 = 7'h23 == io_hh_cnt[6:0] ? myVec_35 : _GEN_74; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_76 = 7'h24 == io_hh_cnt[6:0] ? myVec_36 : _GEN_75; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_77 = 7'h25 == io_hh_cnt[6:0] ? myVec_37 : _GEN_76; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_78 = 7'h26 == io_hh_cnt[6:0] ? myVec_38 : _GEN_77; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_79 = 7'h27 == io_hh_cnt[6:0] ? myVec_39 : _GEN_78; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_80 = 7'h28 == io_hh_cnt[6:0] ? myVec_40 : _GEN_79; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_81 = 7'h29 == io_hh_cnt[6:0] ? myVec_41 : _GEN_80; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_82 = 7'h2a == io_hh_cnt[6:0] ? myVec_42 : _GEN_81; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_83 = 7'h2b == io_hh_cnt[6:0] ? myVec_43 : _GEN_82; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_84 = 7'h2c == io_hh_cnt[6:0] ? myVec_44 : _GEN_83; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_85 = 7'h2d == io_hh_cnt[6:0] ? myVec_45 : _GEN_84; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_86 = 7'h2e == io_hh_cnt[6:0] ? myVec_46 : _GEN_85; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_87 = 7'h2f == io_hh_cnt[6:0] ? myVec_47 : _GEN_86; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_88 = 7'h30 == io_hh_cnt[6:0] ? myVec_48 : _GEN_87; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_89 = 7'h31 == io_hh_cnt[6:0] ? myVec_49 : _GEN_88; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_90 = 7'h32 == io_hh_cnt[6:0] ? myVec_50 : _GEN_89; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_91 = 7'h33 == io_hh_cnt[6:0] ? myVec_51 : _GEN_90; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_92 = 7'h34 == io_hh_cnt[6:0] ? myVec_52 : _GEN_91; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_93 = 7'h35 == io_hh_cnt[6:0] ? myVec_53 : _GEN_92; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_94 = 7'h36 == io_hh_cnt[6:0] ? myVec_54 : _GEN_93; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_95 = 7'h37 == io_hh_cnt[6:0] ? myVec_55 : _GEN_94; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_96 = 7'h38 == io_hh_cnt[6:0] ? myVec_56 : _GEN_95; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_97 = 7'h39 == io_hh_cnt[6:0] ? myVec_57 : _GEN_96; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_98 = 7'h3a == io_hh_cnt[6:0] ? myVec_58 : _GEN_97; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_99 = 7'h3b == io_hh_cnt[6:0] ? myVec_59 : _GEN_98; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_100 = 7'h3c == io_hh_cnt[6:0] ? myVec_60 : _GEN_99; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_101 = 7'h3d == io_hh_cnt[6:0] ? myVec_61 : _GEN_100; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_102 = 7'h3e == io_hh_cnt[6:0] ? myVec_62 : _GEN_101; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_103 = 7'h3f == io_hh_cnt[6:0] ? myVec_63 : _GEN_102; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_104 = 7'h40 == io_hh_cnt[6:0] ? myVec_64 : _GEN_103; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_105 = 7'h41 == io_hh_cnt[6:0] ? myVec_65 : _GEN_104; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_106 = 7'h42 == io_hh_cnt[6:0] ? myVec_66 : _GEN_105; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_107 = 7'h43 == io_hh_cnt[6:0] ? myVec_67 : _GEN_106; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_108 = 7'h44 == io_hh_cnt[6:0] ? myVec_68 : _GEN_107; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_109 = 7'h45 == io_hh_cnt[6:0] ? myVec_69 : _GEN_108; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_110 = 7'h46 == io_hh_cnt[6:0] ? myVec_70 : _GEN_109; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_111 = 7'h47 == io_hh_cnt[6:0] ? myVec_71 : _GEN_110; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_112 = 7'h48 == io_hh_cnt[6:0] ? myVec_72 : _GEN_111; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_113 = 7'h49 == io_hh_cnt[6:0] ? myVec_73 : _GEN_112; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_114 = 7'h4a == io_hh_cnt[6:0] ? myVec_74 : _GEN_113; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_115 = 7'h4b == io_hh_cnt[6:0] ? myVec_75 : _GEN_114; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_116 = 7'h4c == io_hh_cnt[6:0] ? myVec_76 : _GEN_115; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_117 = 7'h4d == io_hh_cnt[6:0] ? myVec_77 : _GEN_116; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_118 = 7'h4e == io_hh_cnt[6:0] ? myVec_78 : _GEN_117; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_119 = 7'h4f == io_hh_cnt[6:0] ? myVec_79 : _GEN_118; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_120 = 7'h50 == io_hh_cnt[6:0] ? myVec_80 : _GEN_119; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_121 = 7'h51 == io_hh_cnt[6:0] ? myVec_81 : _GEN_120; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_122 = 7'h52 == io_hh_cnt[6:0] ? myVec_82 : _GEN_121; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_123 = 7'h53 == io_hh_cnt[6:0] ? myVec_83 : _GEN_122; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_124 = 7'h54 == io_hh_cnt[6:0] ? myVec_84 : _GEN_123; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_125 = 7'h55 == io_hh_cnt[6:0] ? myVec_85 : _GEN_124; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_126 = 7'h56 == io_hh_cnt[6:0] ? myVec_86 : _GEN_125; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_127 = 7'h57 == io_hh_cnt[6:0] ? myVec_87 : _GEN_126; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_128 = 7'h58 == io_hh_cnt[6:0] ? myVec_88 : _GEN_127; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_129 = 7'h59 == io_hh_cnt[6:0] ? myVec_89 : _GEN_128; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_130 = 7'h5a == io_hh_cnt[6:0] ? myVec_90 : _GEN_129; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_131 = 7'h5b == io_hh_cnt[6:0] ? myVec_91 : _GEN_130; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_132 = 7'h5c == io_hh_cnt[6:0] ? myVec_92 : _GEN_131; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_133 = 7'h5d == io_hh_cnt[6:0] ? myVec_93 : _GEN_132; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_134 = 7'h5e == io_hh_cnt[6:0] ? myVec_94 : _GEN_133; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_135 = 7'h5f == io_hh_cnt[6:0] ? myVec_95 : _GEN_134; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_136 = 7'h60 == io_hh_cnt[6:0] ? myVec_96 : _GEN_135; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_137 = 7'h61 == io_hh_cnt[6:0] ? myVec_97 : _GEN_136; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_138 = 7'h62 == io_hh_cnt[6:0] ? myVec_98 : _GEN_137; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_139 = 7'h63 == io_hh_cnt[6:0] ? myVec_99 : _GEN_138; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_140 = 7'h64 == io_hh_cnt[6:0] ? myVec_100 : _GEN_139; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_141 = 7'h65 == io_hh_cnt[6:0] ? myVec_101 : _GEN_140; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_142 = 7'h66 == io_hh_cnt[6:0] ? myVec_102 : _GEN_141; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_143 = 7'h67 == io_hh_cnt[6:0] ? myVec_103 : _GEN_142; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_144 = 7'h68 == io_hh_cnt[6:0] ? myVec_104 : _GEN_143; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_145 = 7'h69 == io_hh_cnt[6:0] ? myVec_105 : _GEN_144; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_146 = 7'h6a == io_hh_cnt[6:0] ? myVec_106 : _GEN_145; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_147 = 7'h6b == io_hh_cnt[6:0] ? myVec_107 : _GEN_146; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_148 = 7'h6c == io_hh_cnt[6:0] ? myVec_108 : _GEN_147; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_149 = 7'h6d == io_hh_cnt[6:0] ? myVec_109 : _GEN_148; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_150 = 7'h6e == io_hh_cnt[6:0] ? myVec_110 : _GEN_149; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_151 = 7'h6f == io_hh_cnt[6:0] ? myVec_111 : _GEN_150; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_152 = 7'h70 == io_hh_cnt[6:0] ? myVec_112 : _GEN_151; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_153 = 7'h71 == io_hh_cnt[6:0] ? myVec_113 : _GEN_152; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_154 = 7'h72 == io_hh_cnt[6:0] ? myVec_114 : _GEN_153; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_155 = 7'h73 == io_hh_cnt[6:0] ? myVec_115 : _GEN_154; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_156 = 7'h74 == io_hh_cnt[6:0] ? myVec_116 : _GEN_155; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_157 = 7'h75 == io_hh_cnt[6:0] ? myVec_117 : _GEN_156; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_158 = 7'h76 == io_hh_cnt[6:0] ? myVec_118 : _GEN_157; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_159 = 7'h77 == io_hh_cnt[6:0] ? myVec_119 : _GEN_158; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_160 = 7'h78 == io_hh_cnt[6:0] ? myVec_120 : _GEN_159; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_161 = 7'h79 == io_hh_cnt[6:0] ? myVec_121 : _GEN_160; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_162 = 7'h7a == io_hh_cnt[6:0] ? myVec_122 : _GEN_161; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_163 = 7'h7b == io_hh_cnt[6:0] ? myVec_123 : _GEN_162; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_164 = 7'h7c == io_hh_cnt[6:0] ? myVec_124 : _GEN_163; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_165 = 7'h7d == io_hh_cnt[6:0] ? myVec_125 : _GEN_164; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_166 = 7'h7e == io_hh_cnt[6:0] ? myVec_126 : _GEN_165; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_167 = 7'h7f == io_hh_cnt[6:0] ? myVec_127 : _GEN_166; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_168 = io_d1_rdy ? _GEN_167 : 32'h0; // @[hh_datapath_chisel.scala 225:26 226:17 228:17]
  wire [31:0] x1_update = io_rst ? 32'h0 : _GEN_168; // @[hh_datapath_chisel.scala 223:17 224:17]
  wire [31:0] d2_update = FP_square_root_newfpu_io_out_s; // @[hh_datapath_chisel.scala 259:15 90:25]
  wire [31:0] tk_update = hqr7_io_out_s; // @[hh_datapath_chisel.scala 268:14 92:25]
  wire [31:0] d5_update = FP_multiplier_10ccs_io_out_s; // @[hh_datapath_chisel.scala 274:14 94:25]
  reg [4063:0] d4_update_reg; // @[hh_datapath_chisel.scala 161:28]
  wire [4095:0] _d4_update_reg_T = {ddot_dout,d4_update_reg}; // @[Cat.scala 31:58]
  wire [31:0] myAxpyVec_1 = axpy_dp_io_out_s_126; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_0 = axpy_dp_io_out_s_127; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_3 = axpy_dp_io_out_s_124; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_2 = axpy_dp_io_out_s_125; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_5 = axpy_dp_io_out_s_122; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_4 = axpy_dp_io_out_s_123; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_7 = axpy_dp_io_out_s_120; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_6 = axpy_dp_io_out_s_121; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [255:0] io_hh_dout_lo_lo_lo_lo = {myAxpyVec_7,myAxpyVec_6,myAxpyVec_5,myAxpyVec_4,myAxpyVec_3,myAxpyVec_2,
    myAxpyVec_1,myAxpyVec_0}; // @[hh_datapath_chisel.scala 286:28]
  wire [31:0] myAxpyVec_9 = axpy_dp_io_out_s_118; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_8 = axpy_dp_io_out_s_119; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_11 = axpy_dp_io_out_s_116; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_10 = axpy_dp_io_out_s_117; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_13 = axpy_dp_io_out_s_114; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_12 = axpy_dp_io_out_s_115; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_15 = axpy_dp_io_out_s_112; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_14 = axpy_dp_io_out_s_113; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [511:0] io_hh_dout_lo_lo_lo = {myAxpyVec_15,myAxpyVec_14,myAxpyVec_13,myAxpyVec_12,myAxpyVec_11,myAxpyVec_10,
    myAxpyVec_9,myAxpyVec_8,io_hh_dout_lo_lo_lo_lo}; // @[hh_datapath_chisel.scala 286:28]
  wire [31:0] myAxpyVec_17 = axpy_dp_io_out_s_110; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_16 = axpy_dp_io_out_s_111; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_19 = axpy_dp_io_out_s_108; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_18 = axpy_dp_io_out_s_109; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_21 = axpy_dp_io_out_s_106; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_20 = axpy_dp_io_out_s_107; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_23 = axpy_dp_io_out_s_104; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_22 = axpy_dp_io_out_s_105; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [255:0] io_hh_dout_lo_lo_hi_lo = {myAxpyVec_23,myAxpyVec_22,myAxpyVec_21,myAxpyVec_20,myAxpyVec_19,myAxpyVec_18,
    myAxpyVec_17,myAxpyVec_16}; // @[hh_datapath_chisel.scala 286:28]
  wire [31:0] myAxpyVec_25 = axpy_dp_io_out_s_102; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_24 = axpy_dp_io_out_s_103; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_27 = axpy_dp_io_out_s_100; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_26 = axpy_dp_io_out_s_101; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_29 = axpy_dp_io_out_s_98; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_28 = axpy_dp_io_out_s_99; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_31 = axpy_dp_io_out_s_96; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_30 = axpy_dp_io_out_s_97; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [1023:0] io_hh_dout_lo_lo = {myAxpyVec_31,myAxpyVec_30,myAxpyVec_29,myAxpyVec_28,myAxpyVec_27,myAxpyVec_26,
    myAxpyVec_25,myAxpyVec_24,io_hh_dout_lo_lo_hi_lo,io_hh_dout_lo_lo_lo}; // @[hh_datapath_chisel.scala 286:28]
  wire [31:0] myAxpyVec_33 = axpy_dp_io_out_s_94; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_32 = axpy_dp_io_out_s_95; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_35 = axpy_dp_io_out_s_92; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_34 = axpy_dp_io_out_s_93; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_37 = axpy_dp_io_out_s_90; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_36 = axpy_dp_io_out_s_91; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_39 = axpy_dp_io_out_s_88; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_38 = axpy_dp_io_out_s_89; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [255:0] io_hh_dout_lo_hi_lo_lo = {myAxpyVec_39,myAxpyVec_38,myAxpyVec_37,myAxpyVec_36,myAxpyVec_35,myAxpyVec_34,
    myAxpyVec_33,myAxpyVec_32}; // @[hh_datapath_chisel.scala 286:28]
  wire [31:0] myAxpyVec_41 = axpy_dp_io_out_s_86; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_40 = axpy_dp_io_out_s_87; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_43 = axpy_dp_io_out_s_84; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_42 = axpy_dp_io_out_s_85; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_45 = axpy_dp_io_out_s_82; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_44 = axpy_dp_io_out_s_83; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_47 = axpy_dp_io_out_s_80; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_46 = axpy_dp_io_out_s_81; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [511:0] io_hh_dout_lo_hi_lo = {myAxpyVec_47,myAxpyVec_46,myAxpyVec_45,myAxpyVec_44,myAxpyVec_43,myAxpyVec_42,
    myAxpyVec_41,myAxpyVec_40,io_hh_dout_lo_hi_lo_lo}; // @[hh_datapath_chisel.scala 286:28]
  wire [31:0] myAxpyVec_49 = axpy_dp_io_out_s_78; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_48 = axpy_dp_io_out_s_79; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_51 = axpy_dp_io_out_s_76; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_50 = axpy_dp_io_out_s_77; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_53 = axpy_dp_io_out_s_74; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_52 = axpy_dp_io_out_s_75; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_55 = axpy_dp_io_out_s_72; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_54 = axpy_dp_io_out_s_73; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [255:0] io_hh_dout_lo_hi_hi_lo = {myAxpyVec_55,myAxpyVec_54,myAxpyVec_53,myAxpyVec_52,myAxpyVec_51,myAxpyVec_50,
    myAxpyVec_49,myAxpyVec_48}; // @[hh_datapath_chisel.scala 286:28]
  wire [31:0] myAxpyVec_57 = axpy_dp_io_out_s_70; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_56 = axpy_dp_io_out_s_71; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_59 = axpy_dp_io_out_s_68; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_58 = axpy_dp_io_out_s_69; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_61 = axpy_dp_io_out_s_66; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_60 = axpy_dp_io_out_s_67; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_63 = axpy_dp_io_out_s_64; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_62 = axpy_dp_io_out_s_65; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [1023:0] io_hh_dout_lo_hi = {myAxpyVec_63,myAxpyVec_62,myAxpyVec_61,myAxpyVec_60,myAxpyVec_59,myAxpyVec_58,
    myAxpyVec_57,myAxpyVec_56,io_hh_dout_lo_hi_hi_lo,io_hh_dout_lo_hi_lo}; // @[hh_datapath_chisel.scala 286:28]
  wire [2047:0] io_hh_dout_lo = {io_hh_dout_lo_hi,io_hh_dout_lo_lo}; // @[hh_datapath_chisel.scala 286:28]
  wire [31:0] myAxpyVec_65 = axpy_dp_io_out_s_62; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_64 = axpy_dp_io_out_s_63; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_67 = axpy_dp_io_out_s_60; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_66 = axpy_dp_io_out_s_61; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_69 = axpy_dp_io_out_s_58; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_68 = axpy_dp_io_out_s_59; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_71 = axpy_dp_io_out_s_56; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_70 = axpy_dp_io_out_s_57; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [255:0] io_hh_dout_hi_lo_lo_lo = {myAxpyVec_71,myAxpyVec_70,myAxpyVec_69,myAxpyVec_68,myAxpyVec_67,myAxpyVec_66,
    myAxpyVec_65,myAxpyVec_64}; // @[hh_datapath_chisel.scala 286:28]
  wire [31:0] myAxpyVec_73 = axpy_dp_io_out_s_54; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_72 = axpy_dp_io_out_s_55; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_75 = axpy_dp_io_out_s_52; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_74 = axpy_dp_io_out_s_53; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_77 = axpy_dp_io_out_s_50; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_76 = axpy_dp_io_out_s_51; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_79 = axpy_dp_io_out_s_48; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_78 = axpy_dp_io_out_s_49; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [511:0] io_hh_dout_hi_lo_lo = {myAxpyVec_79,myAxpyVec_78,myAxpyVec_77,myAxpyVec_76,myAxpyVec_75,myAxpyVec_74,
    myAxpyVec_73,myAxpyVec_72,io_hh_dout_hi_lo_lo_lo}; // @[hh_datapath_chisel.scala 286:28]
  wire [31:0] myAxpyVec_81 = axpy_dp_io_out_s_46; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_80 = axpy_dp_io_out_s_47; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_83 = axpy_dp_io_out_s_44; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_82 = axpy_dp_io_out_s_45; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_85 = axpy_dp_io_out_s_42; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_84 = axpy_dp_io_out_s_43; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_87 = axpy_dp_io_out_s_40; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_86 = axpy_dp_io_out_s_41; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [255:0] io_hh_dout_hi_lo_hi_lo = {myAxpyVec_87,myAxpyVec_86,myAxpyVec_85,myAxpyVec_84,myAxpyVec_83,myAxpyVec_82,
    myAxpyVec_81,myAxpyVec_80}; // @[hh_datapath_chisel.scala 286:28]
  wire [31:0] myAxpyVec_89 = axpy_dp_io_out_s_38; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_88 = axpy_dp_io_out_s_39; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_91 = axpy_dp_io_out_s_36; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_90 = axpy_dp_io_out_s_37; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_93 = axpy_dp_io_out_s_34; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_92 = axpy_dp_io_out_s_35; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_95 = axpy_dp_io_out_s_32; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_94 = axpy_dp_io_out_s_33; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [1023:0] io_hh_dout_hi_lo = {myAxpyVec_95,myAxpyVec_94,myAxpyVec_93,myAxpyVec_92,myAxpyVec_91,myAxpyVec_90,
    myAxpyVec_89,myAxpyVec_88,io_hh_dout_hi_lo_hi_lo,io_hh_dout_hi_lo_lo}; // @[hh_datapath_chisel.scala 286:28]
  wire [31:0] myAxpyVec_97 = axpy_dp_io_out_s_30; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_96 = axpy_dp_io_out_s_31; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_99 = axpy_dp_io_out_s_28; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_98 = axpy_dp_io_out_s_29; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_101 = axpy_dp_io_out_s_26; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_100 = axpy_dp_io_out_s_27; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_103 = axpy_dp_io_out_s_24; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_102 = axpy_dp_io_out_s_25; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [255:0] io_hh_dout_hi_hi_lo_lo = {myAxpyVec_103,myAxpyVec_102,myAxpyVec_101,myAxpyVec_100,myAxpyVec_99,
    myAxpyVec_98,myAxpyVec_97,myAxpyVec_96}; // @[hh_datapath_chisel.scala 286:28]
  wire [31:0] myAxpyVec_105 = axpy_dp_io_out_s_22; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_104 = axpy_dp_io_out_s_23; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_107 = axpy_dp_io_out_s_20; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_106 = axpy_dp_io_out_s_21; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_109 = axpy_dp_io_out_s_18; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_108 = axpy_dp_io_out_s_19; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_111 = axpy_dp_io_out_s_16; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_110 = axpy_dp_io_out_s_17; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [511:0] io_hh_dout_hi_hi_lo = {myAxpyVec_111,myAxpyVec_110,myAxpyVec_109,myAxpyVec_108,myAxpyVec_107,
    myAxpyVec_106,myAxpyVec_105,myAxpyVec_104,io_hh_dout_hi_hi_lo_lo}; // @[hh_datapath_chisel.scala 286:28]
  wire [31:0] myAxpyVec_113 = axpy_dp_io_out_s_14; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_112 = axpy_dp_io_out_s_15; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_115 = axpy_dp_io_out_s_12; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_114 = axpy_dp_io_out_s_13; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_117 = axpy_dp_io_out_s_10; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_116 = axpy_dp_io_out_s_11; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_119 = axpy_dp_io_out_s_8; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_118 = axpy_dp_io_out_s_9; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [255:0] io_hh_dout_hi_hi_hi_lo = {myAxpyVec_119,myAxpyVec_118,myAxpyVec_117,myAxpyVec_116,myAxpyVec_115,
    myAxpyVec_114,myAxpyVec_113,myAxpyVec_112}; // @[hh_datapath_chisel.scala 286:28]
  wire [31:0] myAxpyVec_121 = axpy_dp_io_out_s_6; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_120 = axpy_dp_io_out_s_7; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_123 = axpy_dp_io_out_s_4; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_122 = axpy_dp_io_out_s_5; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_125 = axpy_dp_io_out_s_2; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_124 = axpy_dp_io_out_s_3; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_127 = axpy_dp_io_out_s_0; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [31:0] myAxpyVec_126 = axpy_dp_io_out_s_1; // @[hh_datapath_chisel.scala 282:24 284:36]
  wire [1023:0] io_hh_dout_hi_hi = {myAxpyVec_127,myAxpyVec_126,myAxpyVec_125,myAxpyVec_124,myAxpyVec_123,myAxpyVec_122,
    myAxpyVec_121,myAxpyVec_120,io_hh_dout_hi_hi_hi_lo,io_hh_dout_hi_hi_lo}; // @[hh_datapath_chisel.scala 286:28]
  wire [2047:0] io_hh_dout_hi = {io_hh_dout_hi_hi,io_hh_dout_hi_lo}; // @[hh_datapath_chisel.scala 286:28]
  FP_DDOT_dp FP_DDOT_dp ( // @[hh_datapath_chisel.scala 248:21]
    .clock(FP_DDOT_dp_clock),
    .reset(FP_DDOT_dp_reset),
    .io_in_a_0(FP_DDOT_dp_io_in_a_0),
    .io_in_a_1(FP_DDOT_dp_io_in_a_1),
    .io_in_a_2(FP_DDOT_dp_io_in_a_2),
    .io_in_a_3(FP_DDOT_dp_io_in_a_3),
    .io_in_a_4(FP_DDOT_dp_io_in_a_4),
    .io_in_a_5(FP_DDOT_dp_io_in_a_5),
    .io_in_a_6(FP_DDOT_dp_io_in_a_6),
    .io_in_a_7(FP_DDOT_dp_io_in_a_7),
    .io_in_a_8(FP_DDOT_dp_io_in_a_8),
    .io_in_a_9(FP_DDOT_dp_io_in_a_9),
    .io_in_a_10(FP_DDOT_dp_io_in_a_10),
    .io_in_a_11(FP_DDOT_dp_io_in_a_11),
    .io_in_a_12(FP_DDOT_dp_io_in_a_12),
    .io_in_a_13(FP_DDOT_dp_io_in_a_13),
    .io_in_a_14(FP_DDOT_dp_io_in_a_14),
    .io_in_a_15(FP_DDOT_dp_io_in_a_15),
    .io_in_a_16(FP_DDOT_dp_io_in_a_16),
    .io_in_a_17(FP_DDOT_dp_io_in_a_17),
    .io_in_a_18(FP_DDOT_dp_io_in_a_18),
    .io_in_a_19(FP_DDOT_dp_io_in_a_19),
    .io_in_a_20(FP_DDOT_dp_io_in_a_20),
    .io_in_a_21(FP_DDOT_dp_io_in_a_21),
    .io_in_a_22(FP_DDOT_dp_io_in_a_22),
    .io_in_a_23(FP_DDOT_dp_io_in_a_23),
    .io_in_a_24(FP_DDOT_dp_io_in_a_24),
    .io_in_a_25(FP_DDOT_dp_io_in_a_25),
    .io_in_a_26(FP_DDOT_dp_io_in_a_26),
    .io_in_a_27(FP_DDOT_dp_io_in_a_27),
    .io_in_a_28(FP_DDOT_dp_io_in_a_28),
    .io_in_a_29(FP_DDOT_dp_io_in_a_29),
    .io_in_a_30(FP_DDOT_dp_io_in_a_30),
    .io_in_a_31(FP_DDOT_dp_io_in_a_31),
    .io_in_a_32(FP_DDOT_dp_io_in_a_32),
    .io_in_a_33(FP_DDOT_dp_io_in_a_33),
    .io_in_a_34(FP_DDOT_dp_io_in_a_34),
    .io_in_a_35(FP_DDOT_dp_io_in_a_35),
    .io_in_a_36(FP_DDOT_dp_io_in_a_36),
    .io_in_a_37(FP_DDOT_dp_io_in_a_37),
    .io_in_a_38(FP_DDOT_dp_io_in_a_38),
    .io_in_a_39(FP_DDOT_dp_io_in_a_39),
    .io_in_a_40(FP_DDOT_dp_io_in_a_40),
    .io_in_a_41(FP_DDOT_dp_io_in_a_41),
    .io_in_a_42(FP_DDOT_dp_io_in_a_42),
    .io_in_a_43(FP_DDOT_dp_io_in_a_43),
    .io_in_a_44(FP_DDOT_dp_io_in_a_44),
    .io_in_a_45(FP_DDOT_dp_io_in_a_45),
    .io_in_a_46(FP_DDOT_dp_io_in_a_46),
    .io_in_a_47(FP_DDOT_dp_io_in_a_47),
    .io_in_a_48(FP_DDOT_dp_io_in_a_48),
    .io_in_a_49(FP_DDOT_dp_io_in_a_49),
    .io_in_a_50(FP_DDOT_dp_io_in_a_50),
    .io_in_a_51(FP_DDOT_dp_io_in_a_51),
    .io_in_a_52(FP_DDOT_dp_io_in_a_52),
    .io_in_a_53(FP_DDOT_dp_io_in_a_53),
    .io_in_a_54(FP_DDOT_dp_io_in_a_54),
    .io_in_a_55(FP_DDOT_dp_io_in_a_55),
    .io_in_a_56(FP_DDOT_dp_io_in_a_56),
    .io_in_a_57(FP_DDOT_dp_io_in_a_57),
    .io_in_a_58(FP_DDOT_dp_io_in_a_58),
    .io_in_a_59(FP_DDOT_dp_io_in_a_59),
    .io_in_a_60(FP_DDOT_dp_io_in_a_60),
    .io_in_a_61(FP_DDOT_dp_io_in_a_61),
    .io_in_a_62(FP_DDOT_dp_io_in_a_62),
    .io_in_a_63(FP_DDOT_dp_io_in_a_63),
    .io_in_a_64(FP_DDOT_dp_io_in_a_64),
    .io_in_a_65(FP_DDOT_dp_io_in_a_65),
    .io_in_a_66(FP_DDOT_dp_io_in_a_66),
    .io_in_a_67(FP_DDOT_dp_io_in_a_67),
    .io_in_a_68(FP_DDOT_dp_io_in_a_68),
    .io_in_a_69(FP_DDOT_dp_io_in_a_69),
    .io_in_a_70(FP_DDOT_dp_io_in_a_70),
    .io_in_a_71(FP_DDOT_dp_io_in_a_71),
    .io_in_a_72(FP_DDOT_dp_io_in_a_72),
    .io_in_a_73(FP_DDOT_dp_io_in_a_73),
    .io_in_a_74(FP_DDOT_dp_io_in_a_74),
    .io_in_a_75(FP_DDOT_dp_io_in_a_75),
    .io_in_a_76(FP_DDOT_dp_io_in_a_76),
    .io_in_a_77(FP_DDOT_dp_io_in_a_77),
    .io_in_a_78(FP_DDOT_dp_io_in_a_78),
    .io_in_a_79(FP_DDOT_dp_io_in_a_79),
    .io_in_a_80(FP_DDOT_dp_io_in_a_80),
    .io_in_a_81(FP_DDOT_dp_io_in_a_81),
    .io_in_a_82(FP_DDOT_dp_io_in_a_82),
    .io_in_a_83(FP_DDOT_dp_io_in_a_83),
    .io_in_a_84(FP_DDOT_dp_io_in_a_84),
    .io_in_a_85(FP_DDOT_dp_io_in_a_85),
    .io_in_a_86(FP_DDOT_dp_io_in_a_86),
    .io_in_a_87(FP_DDOT_dp_io_in_a_87),
    .io_in_a_88(FP_DDOT_dp_io_in_a_88),
    .io_in_a_89(FP_DDOT_dp_io_in_a_89),
    .io_in_a_90(FP_DDOT_dp_io_in_a_90),
    .io_in_a_91(FP_DDOT_dp_io_in_a_91),
    .io_in_a_92(FP_DDOT_dp_io_in_a_92),
    .io_in_a_93(FP_DDOT_dp_io_in_a_93),
    .io_in_a_94(FP_DDOT_dp_io_in_a_94),
    .io_in_a_95(FP_DDOT_dp_io_in_a_95),
    .io_in_a_96(FP_DDOT_dp_io_in_a_96),
    .io_in_a_97(FP_DDOT_dp_io_in_a_97),
    .io_in_a_98(FP_DDOT_dp_io_in_a_98),
    .io_in_a_99(FP_DDOT_dp_io_in_a_99),
    .io_in_a_100(FP_DDOT_dp_io_in_a_100),
    .io_in_a_101(FP_DDOT_dp_io_in_a_101),
    .io_in_a_102(FP_DDOT_dp_io_in_a_102),
    .io_in_a_103(FP_DDOT_dp_io_in_a_103),
    .io_in_a_104(FP_DDOT_dp_io_in_a_104),
    .io_in_a_105(FP_DDOT_dp_io_in_a_105),
    .io_in_a_106(FP_DDOT_dp_io_in_a_106),
    .io_in_a_107(FP_DDOT_dp_io_in_a_107),
    .io_in_a_108(FP_DDOT_dp_io_in_a_108),
    .io_in_a_109(FP_DDOT_dp_io_in_a_109),
    .io_in_a_110(FP_DDOT_dp_io_in_a_110),
    .io_in_a_111(FP_DDOT_dp_io_in_a_111),
    .io_in_a_112(FP_DDOT_dp_io_in_a_112),
    .io_in_a_113(FP_DDOT_dp_io_in_a_113),
    .io_in_a_114(FP_DDOT_dp_io_in_a_114),
    .io_in_a_115(FP_DDOT_dp_io_in_a_115),
    .io_in_a_116(FP_DDOT_dp_io_in_a_116),
    .io_in_a_117(FP_DDOT_dp_io_in_a_117),
    .io_in_a_118(FP_DDOT_dp_io_in_a_118),
    .io_in_a_119(FP_DDOT_dp_io_in_a_119),
    .io_in_a_120(FP_DDOT_dp_io_in_a_120),
    .io_in_a_121(FP_DDOT_dp_io_in_a_121),
    .io_in_a_122(FP_DDOT_dp_io_in_a_122),
    .io_in_a_123(FP_DDOT_dp_io_in_a_123),
    .io_in_a_124(FP_DDOT_dp_io_in_a_124),
    .io_in_a_125(FP_DDOT_dp_io_in_a_125),
    .io_in_a_126(FP_DDOT_dp_io_in_a_126),
    .io_in_a_127(FP_DDOT_dp_io_in_a_127),
    .io_in_b_0(FP_DDOT_dp_io_in_b_0),
    .io_in_b_1(FP_DDOT_dp_io_in_b_1),
    .io_in_b_2(FP_DDOT_dp_io_in_b_2),
    .io_in_b_3(FP_DDOT_dp_io_in_b_3),
    .io_in_b_4(FP_DDOT_dp_io_in_b_4),
    .io_in_b_5(FP_DDOT_dp_io_in_b_5),
    .io_in_b_6(FP_DDOT_dp_io_in_b_6),
    .io_in_b_7(FP_DDOT_dp_io_in_b_7),
    .io_in_b_8(FP_DDOT_dp_io_in_b_8),
    .io_in_b_9(FP_DDOT_dp_io_in_b_9),
    .io_in_b_10(FP_DDOT_dp_io_in_b_10),
    .io_in_b_11(FP_DDOT_dp_io_in_b_11),
    .io_in_b_12(FP_DDOT_dp_io_in_b_12),
    .io_in_b_13(FP_DDOT_dp_io_in_b_13),
    .io_in_b_14(FP_DDOT_dp_io_in_b_14),
    .io_in_b_15(FP_DDOT_dp_io_in_b_15),
    .io_in_b_16(FP_DDOT_dp_io_in_b_16),
    .io_in_b_17(FP_DDOT_dp_io_in_b_17),
    .io_in_b_18(FP_DDOT_dp_io_in_b_18),
    .io_in_b_19(FP_DDOT_dp_io_in_b_19),
    .io_in_b_20(FP_DDOT_dp_io_in_b_20),
    .io_in_b_21(FP_DDOT_dp_io_in_b_21),
    .io_in_b_22(FP_DDOT_dp_io_in_b_22),
    .io_in_b_23(FP_DDOT_dp_io_in_b_23),
    .io_in_b_24(FP_DDOT_dp_io_in_b_24),
    .io_in_b_25(FP_DDOT_dp_io_in_b_25),
    .io_in_b_26(FP_DDOT_dp_io_in_b_26),
    .io_in_b_27(FP_DDOT_dp_io_in_b_27),
    .io_in_b_28(FP_DDOT_dp_io_in_b_28),
    .io_in_b_29(FP_DDOT_dp_io_in_b_29),
    .io_in_b_30(FP_DDOT_dp_io_in_b_30),
    .io_in_b_31(FP_DDOT_dp_io_in_b_31),
    .io_in_b_32(FP_DDOT_dp_io_in_b_32),
    .io_in_b_33(FP_DDOT_dp_io_in_b_33),
    .io_in_b_34(FP_DDOT_dp_io_in_b_34),
    .io_in_b_35(FP_DDOT_dp_io_in_b_35),
    .io_in_b_36(FP_DDOT_dp_io_in_b_36),
    .io_in_b_37(FP_DDOT_dp_io_in_b_37),
    .io_in_b_38(FP_DDOT_dp_io_in_b_38),
    .io_in_b_39(FP_DDOT_dp_io_in_b_39),
    .io_in_b_40(FP_DDOT_dp_io_in_b_40),
    .io_in_b_41(FP_DDOT_dp_io_in_b_41),
    .io_in_b_42(FP_DDOT_dp_io_in_b_42),
    .io_in_b_43(FP_DDOT_dp_io_in_b_43),
    .io_in_b_44(FP_DDOT_dp_io_in_b_44),
    .io_in_b_45(FP_DDOT_dp_io_in_b_45),
    .io_in_b_46(FP_DDOT_dp_io_in_b_46),
    .io_in_b_47(FP_DDOT_dp_io_in_b_47),
    .io_in_b_48(FP_DDOT_dp_io_in_b_48),
    .io_in_b_49(FP_DDOT_dp_io_in_b_49),
    .io_in_b_50(FP_DDOT_dp_io_in_b_50),
    .io_in_b_51(FP_DDOT_dp_io_in_b_51),
    .io_in_b_52(FP_DDOT_dp_io_in_b_52),
    .io_in_b_53(FP_DDOT_dp_io_in_b_53),
    .io_in_b_54(FP_DDOT_dp_io_in_b_54),
    .io_in_b_55(FP_DDOT_dp_io_in_b_55),
    .io_in_b_56(FP_DDOT_dp_io_in_b_56),
    .io_in_b_57(FP_DDOT_dp_io_in_b_57),
    .io_in_b_58(FP_DDOT_dp_io_in_b_58),
    .io_in_b_59(FP_DDOT_dp_io_in_b_59),
    .io_in_b_60(FP_DDOT_dp_io_in_b_60),
    .io_in_b_61(FP_DDOT_dp_io_in_b_61),
    .io_in_b_62(FP_DDOT_dp_io_in_b_62),
    .io_in_b_63(FP_DDOT_dp_io_in_b_63),
    .io_in_b_64(FP_DDOT_dp_io_in_b_64),
    .io_in_b_65(FP_DDOT_dp_io_in_b_65),
    .io_in_b_66(FP_DDOT_dp_io_in_b_66),
    .io_in_b_67(FP_DDOT_dp_io_in_b_67),
    .io_in_b_68(FP_DDOT_dp_io_in_b_68),
    .io_in_b_69(FP_DDOT_dp_io_in_b_69),
    .io_in_b_70(FP_DDOT_dp_io_in_b_70),
    .io_in_b_71(FP_DDOT_dp_io_in_b_71),
    .io_in_b_72(FP_DDOT_dp_io_in_b_72),
    .io_in_b_73(FP_DDOT_dp_io_in_b_73),
    .io_in_b_74(FP_DDOT_dp_io_in_b_74),
    .io_in_b_75(FP_DDOT_dp_io_in_b_75),
    .io_in_b_76(FP_DDOT_dp_io_in_b_76),
    .io_in_b_77(FP_DDOT_dp_io_in_b_77),
    .io_in_b_78(FP_DDOT_dp_io_in_b_78),
    .io_in_b_79(FP_DDOT_dp_io_in_b_79),
    .io_in_b_80(FP_DDOT_dp_io_in_b_80),
    .io_in_b_81(FP_DDOT_dp_io_in_b_81),
    .io_in_b_82(FP_DDOT_dp_io_in_b_82),
    .io_in_b_83(FP_DDOT_dp_io_in_b_83),
    .io_in_b_84(FP_DDOT_dp_io_in_b_84),
    .io_in_b_85(FP_DDOT_dp_io_in_b_85),
    .io_in_b_86(FP_DDOT_dp_io_in_b_86),
    .io_in_b_87(FP_DDOT_dp_io_in_b_87),
    .io_in_b_88(FP_DDOT_dp_io_in_b_88),
    .io_in_b_89(FP_DDOT_dp_io_in_b_89),
    .io_in_b_90(FP_DDOT_dp_io_in_b_90),
    .io_in_b_91(FP_DDOT_dp_io_in_b_91),
    .io_in_b_92(FP_DDOT_dp_io_in_b_92),
    .io_in_b_93(FP_DDOT_dp_io_in_b_93),
    .io_in_b_94(FP_DDOT_dp_io_in_b_94),
    .io_in_b_95(FP_DDOT_dp_io_in_b_95),
    .io_in_b_96(FP_DDOT_dp_io_in_b_96),
    .io_in_b_97(FP_DDOT_dp_io_in_b_97),
    .io_in_b_98(FP_DDOT_dp_io_in_b_98),
    .io_in_b_99(FP_DDOT_dp_io_in_b_99),
    .io_in_b_100(FP_DDOT_dp_io_in_b_100),
    .io_in_b_101(FP_DDOT_dp_io_in_b_101),
    .io_in_b_102(FP_DDOT_dp_io_in_b_102),
    .io_in_b_103(FP_DDOT_dp_io_in_b_103),
    .io_in_b_104(FP_DDOT_dp_io_in_b_104),
    .io_in_b_105(FP_DDOT_dp_io_in_b_105),
    .io_in_b_106(FP_DDOT_dp_io_in_b_106),
    .io_in_b_107(FP_DDOT_dp_io_in_b_107),
    .io_in_b_108(FP_DDOT_dp_io_in_b_108),
    .io_in_b_109(FP_DDOT_dp_io_in_b_109),
    .io_in_b_110(FP_DDOT_dp_io_in_b_110),
    .io_in_b_111(FP_DDOT_dp_io_in_b_111),
    .io_in_b_112(FP_DDOT_dp_io_in_b_112),
    .io_in_b_113(FP_DDOT_dp_io_in_b_113),
    .io_in_b_114(FP_DDOT_dp_io_in_b_114),
    .io_in_b_115(FP_DDOT_dp_io_in_b_115),
    .io_in_b_116(FP_DDOT_dp_io_in_b_116),
    .io_in_b_117(FP_DDOT_dp_io_in_b_117),
    .io_in_b_118(FP_DDOT_dp_io_in_b_118),
    .io_in_b_119(FP_DDOT_dp_io_in_b_119),
    .io_in_b_120(FP_DDOT_dp_io_in_b_120),
    .io_in_b_121(FP_DDOT_dp_io_in_b_121),
    .io_in_b_122(FP_DDOT_dp_io_in_b_122),
    .io_in_b_123(FP_DDOT_dp_io_in_b_123),
    .io_in_b_124(FP_DDOT_dp_io_in_b_124),
    .io_in_b_125(FP_DDOT_dp_io_in_b_125),
    .io_in_b_126(FP_DDOT_dp_io_in_b_126),
    .io_in_b_127(FP_DDOT_dp_io_in_b_127),
    .io_out_s(FP_DDOT_dp_io_out_s)
  );
  FP_square_root_newfpu FP_square_root_newfpu ( // @[hh_datapath_chisel.scala 256:22]
    .clock(FP_square_root_newfpu_clock),
    .reset(FP_square_root_newfpu_reset),
    .io_in_a(FP_square_root_newfpu_io_in_a),
    .io_out_s(FP_square_root_newfpu_io_out_s)
  );
  hqr5 hqr5 ( // @[hh_datapath_chisel.scala 261:20]
    .clock(hqr5_clock),
    .reset(hqr5_reset),
    .io_in_a(hqr5_io_in_a),
    .io_in_b(hqr5_io_in_b),
    .io_out_s(hqr5_io_out_s)
  );
  hqr7 hqr7 ( // @[hh_datapath_chisel.scala 266:20]
    .clock(hqr7_clock),
    .reset(hqr7_reset),
    .io_in_a(hqr7_io_in_a),
    .io_out_s(hqr7_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs ( // @[hh_datapath_chisel.scala 270:21]
    .clock(FP_multiplier_10ccs_clock),
    .reset(FP_multiplier_10ccs_reset),
    .io_in_a(FP_multiplier_10ccs_io_in_a),
    .io_in_b(FP_multiplier_10ccs_io_in_b),
    .io_out_s(FP_multiplier_10ccs_io_out_s)
  );
  axpy_dp axpy_dp ( // @[hh_datapath_chisel.scala 276:20]
    .clock(axpy_dp_clock),
    .reset(axpy_dp_reset),
    .io_in_a(axpy_dp_io_in_a),
    .io_in_b_0(axpy_dp_io_in_b_0),
    .io_in_b_1(axpy_dp_io_in_b_1),
    .io_in_b_2(axpy_dp_io_in_b_2),
    .io_in_b_3(axpy_dp_io_in_b_3),
    .io_in_b_4(axpy_dp_io_in_b_4),
    .io_in_b_5(axpy_dp_io_in_b_5),
    .io_in_b_6(axpy_dp_io_in_b_6),
    .io_in_b_7(axpy_dp_io_in_b_7),
    .io_in_b_8(axpy_dp_io_in_b_8),
    .io_in_b_9(axpy_dp_io_in_b_9),
    .io_in_b_10(axpy_dp_io_in_b_10),
    .io_in_b_11(axpy_dp_io_in_b_11),
    .io_in_b_12(axpy_dp_io_in_b_12),
    .io_in_b_13(axpy_dp_io_in_b_13),
    .io_in_b_14(axpy_dp_io_in_b_14),
    .io_in_b_15(axpy_dp_io_in_b_15),
    .io_in_b_16(axpy_dp_io_in_b_16),
    .io_in_b_17(axpy_dp_io_in_b_17),
    .io_in_b_18(axpy_dp_io_in_b_18),
    .io_in_b_19(axpy_dp_io_in_b_19),
    .io_in_b_20(axpy_dp_io_in_b_20),
    .io_in_b_21(axpy_dp_io_in_b_21),
    .io_in_b_22(axpy_dp_io_in_b_22),
    .io_in_b_23(axpy_dp_io_in_b_23),
    .io_in_b_24(axpy_dp_io_in_b_24),
    .io_in_b_25(axpy_dp_io_in_b_25),
    .io_in_b_26(axpy_dp_io_in_b_26),
    .io_in_b_27(axpy_dp_io_in_b_27),
    .io_in_b_28(axpy_dp_io_in_b_28),
    .io_in_b_29(axpy_dp_io_in_b_29),
    .io_in_b_30(axpy_dp_io_in_b_30),
    .io_in_b_31(axpy_dp_io_in_b_31),
    .io_in_b_32(axpy_dp_io_in_b_32),
    .io_in_b_33(axpy_dp_io_in_b_33),
    .io_in_b_34(axpy_dp_io_in_b_34),
    .io_in_b_35(axpy_dp_io_in_b_35),
    .io_in_b_36(axpy_dp_io_in_b_36),
    .io_in_b_37(axpy_dp_io_in_b_37),
    .io_in_b_38(axpy_dp_io_in_b_38),
    .io_in_b_39(axpy_dp_io_in_b_39),
    .io_in_b_40(axpy_dp_io_in_b_40),
    .io_in_b_41(axpy_dp_io_in_b_41),
    .io_in_b_42(axpy_dp_io_in_b_42),
    .io_in_b_43(axpy_dp_io_in_b_43),
    .io_in_b_44(axpy_dp_io_in_b_44),
    .io_in_b_45(axpy_dp_io_in_b_45),
    .io_in_b_46(axpy_dp_io_in_b_46),
    .io_in_b_47(axpy_dp_io_in_b_47),
    .io_in_b_48(axpy_dp_io_in_b_48),
    .io_in_b_49(axpy_dp_io_in_b_49),
    .io_in_b_50(axpy_dp_io_in_b_50),
    .io_in_b_51(axpy_dp_io_in_b_51),
    .io_in_b_52(axpy_dp_io_in_b_52),
    .io_in_b_53(axpy_dp_io_in_b_53),
    .io_in_b_54(axpy_dp_io_in_b_54),
    .io_in_b_55(axpy_dp_io_in_b_55),
    .io_in_b_56(axpy_dp_io_in_b_56),
    .io_in_b_57(axpy_dp_io_in_b_57),
    .io_in_b_58(axpy_dp_io_in_b_58),
    .io_in_b_59(axpy_dp_io_in_b_59),
    .io_in_b_60(axpy_dp_io_in_b_60),
    .io_in_b_61(axpy_dp_io_in_b_61),
    .io_in_b_62(axpy_dp_io_in_b_62),
    .io_in_b_63(axpy_dp_io_in_b_63),
    .io_in_b_64(axpy_dp_io_in_b_64),
    .io_in_b_65(axpy_dp_io_in_b_65),
    .io_in_b_66(axpy_dp_io_in_b_66),
    .io_in_b_67(axpy_dp_io_in_b_67),
    .io_in_b_68(axpy_dp_io_in_b_68),
    .io_in_b_69(axpy_dp_io_in_b_69),
    .io_in_b_70(axpy_dp_io_in_b_70),
    .io_in_b_71(axpy_dp_io_in_b_71),
    .io_in_b_72(axpy_dp_io_in_b_72),
    .io_in_b_73(axpy_dp_io_in_b_73),
    .io_in_b_74(axpy_dp_io_in_b_74),
    .io_in_b_75(axpy_dp_io_in_b_75),
    .io_in_b_76(axpy_dp_io_in_b_76),
    .io_in_b_77(axpy_dp_io_in_b_77),
    .io_in_b_78(axpy_dp_io_in_b_78),
    .io_in_b_79(axpy_dp_io_in_b_79),
    .io_in_b_80(axpy_dp_io_in_b_80),
    .io_in_b_81(axpy_dp_io_in_b_81),
    .io_in_b_82(axpy_dp_io_in_b_82),
    .io_in_b_83(axpy_dp_io_in_b_83),
    .io_in_b_84(axpy_dp_io_in_b_84),
    .io_in_b_85(axpy_dp_io_in_b_85),
    .io_in_b_86(axpy_dp_io_in_b_86),
    .io_in_b_87(axpy_dp_io_in_b_87),
    .io_in_b_88(axpy_dp_io_in_b_88),
    .io_in_b_89(axpy_dp_io_in_b_89),
    .io_in_b_90(axpy_dp_io_in_b_90),
    .io_in_b_91(axpy_dp_io_in_b_91),
    .io_in_b_92(axpy_dp_io_in_b_92),
    .io_in_b_93(axpy_dp_io_in_b_93),
    .io_in_b_94(axpy_dp_io_in_b_94),
    .io_in_b_95(axpy_dp_io_in_b_95),
    .io_in_b_96(axpy_dp_io_in_b_96),
    .io_in_b_97(axpy_dp_io_in_b_97),
    .io_in_b_98(axpy_dp_io_in_b_98),
    .io_in_b_99(axpy_dp_io_in_b_99),
    .io_in_b_100(axpy_dp_io_in_b_100),
    .io_in_b_101(axpy_dp_io_in_b_101),
    .io_in_b_102(axpy_dp_io_in_b_102),
    .io_in_b_103(axpy_dp_io_in_b_103),
    .io_in_b_104(axpy_dp_io_in_b_104),
    .io_in_b_105(axpy_dp_io_in_b_105),
    .io_in_b_106(axpy_dp_io_in_b_106),
    .io_in_b_107(axpy_dp_io_in_b_107),
    .io_in_b_108(axpy_dp_io_in_b_108),
    .io_in_b_109(axpy_dp_io_in_b_109),
    .io_in_b_110(axpy_dp_io_in_b_110),
    .io_in_b_111(axpy_dp_io_in_b_111),
    .io_in_b_112(axpy_dp_io_in_b_112),
    .io_in_b_113(axpy_dp_io_in_b_113),
    .io_in_b_114(axpy_dp_io_in_b_114),
    .io_in_b_115(axpy_dp_io_in_b_115),
    .io_in_b_116(axpy_dp_io_in_b_116),
    .io_in_b_117(axpy_dp_io_in_b_117),
    .io_in_b_118(axpy_dp_io_in_b_118),
    .io_in_b_119(axpy_dp_io_in_b_119),
    .io_in_b_120(axpy_dp_io_in_b_120),
    .io_in_b_121(axpy_dp_io_in_b_121),
    .io_in_b_122(axpy_dp_io_in_b_122),
    .io_in_b_123(axpy_dp_io_in_b_123),
    .io_in_b_124(axpy_dp_io_in_b_124),
    .io_in_b_125(axpy_dp_io_in_b_125),
    .io_in_b_126(axpy_dp_io_in_b_126),
    .io_in_b_127(axpy_dp_io_in_b_127),
    .io_in_c_0(axpy_dp_io_in_c_0),
    .io_in_c_1(axpy_dp_io_in_c_1),
    .io_in_c_2(axpy_dp_io_in_c_2),
    .io_in_c_3(axpy_dp_io_in_c_3),
    .io_in_c_4(axpy_dp_io_in_c_4),
    .io_in_c_5(axpy_dp_io_in_c_5),
    .io_in_c_6(axpy_dp_io_in_c_6),
    .io_in_c_7(axpy_dp_io_in_c_7),
    .io_in_c_8(axpy_dp_io_in_c_8),
    .io_in_c_9(axpy_dp_io_in_c_9),
    .io_in_c_10(axpy_dp_io_in_c_10),
    .io_in_c_11(axpy_dp_io_in_c_11),
    .io_in_c_12(axpy_dp_io_in_c_12),
    .io_in_c_13(axpy_dp_io_in_c_13),
    .io_in_c_14(axpy_dp_io_in_c_14),
    .io_in_c_15(axpy_dp_io_in_c_15),
    .io_in_c_16(axpy_dp_io_in_c_16),
    .io_in_c_17(axpy_dp_io_in_c_17),
    .io_in_c_18(axpy_dp_io_in_c_18),
    .io_in_c_19(axpy_dp_io_in_c_19),
    .io_in_c_20(axpy_dp_io_in_c_20),
    .io_in_c_21(axpy_dp_io_in_c_21),
    .io_in_c_22(axpy_dp_io_in_c_22),
    .io_in_c_23(axpy_dp_io_in_c_23),
    .io_in_c_24(axpy_dp_io_in_c_24),
    .io_in_c_25(axpy_dp_io_in_c_25),
    .io_in_c_26(axpy_dp_io_in_c_26),
    .io_in_c_27(axpy_dp_io_in_c_27),
    .io_in_c_28(axpy_dp_io_in_c_28),
    .io_in_c_29(axpy_dp_io_in_c_29),
    .io_in_c_30(axpy_dp_io_in_c_30),
    .io_in_c_31(axpy_dp_io_in_c_31),
    .io_in_c_32(axpy_dp_io_in_c_32),
    .io_in_c_33(axpy_dp_io_in_c_33),
    .io_in_c_34(axpy_dp_io_in_c_34),
    .io_in_c_35(axpy_dp_io_in_c_35),
    .io_in_c_36(axpy_dp_io_in_c_36),
    .io_in_c_37(axpy_dp_io_in_c_37),
    .io_in_c_38(axpy_dp_io_in_c_38),
    .io_in_c_39(axpy_dp_io_in_c_39),
    .io_in_c_40(axpy_dp_io_in_c_40),
    .io_in_c_41(axpy_dp_io_in_c_41),
    .io_in_c_42(axpy_dp_io_in_c_42),
    .io_in_c_43(axpy_dp_io_in_c_43),
    .io_in_c_44(axpy_dp_io_in_c_44),
    .io_in_c_45(axpy_dp_io_in_c_45),
    .io_in_c_46(axpy_dp_io_in_c_46),
    .io_in_c_47(axpy_dp_io_in_c_47),
    .io_in_c_48(axpy_dp_io_in_c_48),
    .io_in_c_49(axpy_dp_io_in_c_49),
    .io_in_c_50(axpy_dp_io_in_c_50),
    .io_in_c_51(axpy_dp_io_in_c_51),
    .io_in_c_52(axpy_dp_io_in_c_52),
    .io_in_c_53(axpy_dp_io_in_c_53),
    .io_in_c_54(axpy_dp_io_in_c_54),
    .io_in_c_55(axpy_dp_io_in_c_55),
    .io_in_c_56(axpy_dp_io_in_c_56),
    .io_in_c_57(axpy_dp_io_in_c_57),
    .io_in_c_58(axpy_dp_io_in_c_58),
    .io_in_c_59(axpy_dp_io_in_c_59),
    .io_in_c_60(axpy_dp_io_in_c_60),
    .io_in_c_61(axpy_dp_io_in_c_61),
    .io_in_c_62(axpy_dp_io_in_c_62),
    .io_in_c_63(axpy_dp_io_in_c_63),
    .io_in_c_64(axpy_dp_io_in_c_64),
    .io_in_c_65(axpy_dp_io_in_c_65),
    .io_in_c_66(axpy_dp_io_in_c_66),
    .io_in_c_67(axpy_dp_io_in_c_67),
    .io_in_c_68(axpy_dp_io_in_c_68),
    .io_in_c_69(axpy_dp_io_in_c_69),
    .io_in_c_70(axpy_dp_io_in_c_70),
    .io_in_c_71(axpy_dp_io_in_c_71),
    .io_in_c_72(axpy_dp_io_in_c_72),
    .io_in_c_73(axpy_dp_io_in_c_73),
    .io_in_c_74(axpy_dp_io_in_c_74),
    .io_in_c_75(axpy_dp_io_in_c_75),
    .io_in_c_76(axpy_dp_io_in_c_76),
    .io_in_c_77(axpy_dp_io_in_c_77),
    .io_in_c_78(axpy_dp_io_in_c_78),
    .io_in_c_79(axpy_dp_io_in_c_79),
    .io_in_c_80(axpy_dp_io_in_c_80),
    .io_in_c_81(axpy_dp_io_in_c_81),
    .io_in_c_82(axpy_dp_io_in_c_82),
    .io_in_c_83(axpy_dp_io_in_c_83),
    .io_in_c_84(axpy_dp_io_in_c_84),
    .io_in_c_85(axpy_dp_io_in_c_85),
    .io_in_c_86(axpy_dp_io_in_c_86),
    .io_in_c_87(axpy_dp_io_in_c_87),
    .io_in_c_88(axpy_dp_io_in_c_88),
    .io_in_c_89(axpy_dp_io_in_c_89),
    .io_in_c_90(axpy_dp_io_in_c_90),
    .io_in_c_91(axpy_dp_io_in_c_91),
    .io_in_c_92(axpy_dp_io_in_c_92),
    .io_in_c_93(axpy_dp_io_in_c_93),
    .io_in_c_94(axpy_dp_io_in_c_94),
    .io_in_c_95(axpy_dp_io_in_c_95),
    .io_in_c_96(axpy_dp_io_in_c_96),
    .io_in_c_97(axpy_dp_io_in_c_97),
    .io_in_c_98(axpy_dp_io_in_c_98),
    .io_in_c_99(axpy_dp_io_in_c_99),
    .io_in_c_100(axpy_dp_io_in_c_100),
    .io_in_c_101(axpy_dp_io_in_c_101),
    .io_in_c_102(axpy_dp_io_in_c_102),
    .io_in_c_103(axpy_dp_io_in_c_103),
    .io_in_c_104(axpy_dp_io_in_c_104),
    .io_in_c_105(axpy_dp_io_in_c_105),
    .io_in_c_106(axpy_dp_io_in_c_106),
    .io_in_c_107(axpy_dp_io_in_c_107),
    .io_in_c_108(axpy_dp_io_in_c_108),
    .io_in_c_109(axpy_dp_io_in_c_109),
    .io_in_c_110(axpy_dp_io_in_c_110),
    .io_in_c_111(axpy_dp_io_in_c_111),
    .io_in_c_112(axpy_dp_io_in_c_112),
    .io_in_c_113(axpy_dp_io_in_c_113),
    .io_in_c_114(axpy_dp_io_in_c_114),
    .io_in_c_115(axpy_dp_io_in_c_115),
    .io_in_c_116(axpy_dp_io_in_c_116),
    .io_in_c_117(axpy_dp_io_in_c_117),
    .io_in_c_118(axpy_dp_io_in_c_118),
    .io_in_c_119(axpy_dp_io_in_c_119),
    .io_in_c_120(axpy_dp_io_in_c_120),
    .io_in_c_121(axpy_dp_io_in_c_121),
    .io_in_c_122(axpy_dp_io_in_c_122),
    .io_in_c_123(axpy_dp_io_in_c_123),
    .io_in_c_124(axpy_dp_io_in_c_124),
    .io_in_c_125(axpy_dp_io_in_c_125),
    .io_in_c_126(axpy_dp_io_in_c_126),
    .io_in_c_127(axpy_dp_io_in_c_127),
    .io_out_s_0(axpy_dp_io_out_s_0),
    .io_out_s_1(axpy_dp_io_out_s_1),
    .io_out_s_2(axpy_dp_io_out_s_2),
    .io_out_s_3(axpy_dp_io_out_s_3),
    .io_out_s_4(axpy_dp_io_out_s_4),
    .io_out_s_5(axpy_dp_io_out_s_5),
    .io_out_s_6(axpy_dp_io_out_s_6),
    .io_out_s_7(axpy_dp_io_out_s_7),
    .io_out_s_8(axpy_dp_io_out_s_8),
    .io_out_s_9(axpy_dp_io_out_s_9),
    .io_out_s_10(axpy_dp_io_out_s_10),
    .io_out_s_11(axpy_dp_io_out_s_11),
    .io_out_s_12(axpy_dp_io_out_s_12),
    .io_out_s_13(axpy_dp_io_out_s_13),
    .io_out_s_14(axpy_dp_io_out_s_14),
    .io_out_s_15(axpy_dp_io_out_s_15),
    .io_out_s_16(axpy_dp_io_out_s_16),
    .io_out_s_17(axpy_dp_io_out_s_17),
    .io_out_s_18(axpy_dp_io_out_s_18),
    .io_out_s_19(axpy_dp_io_out_s_19),
    .io_out_s_20(axpy_dp_io_out_s_20),
    .io_out_s_21(axpy_dp_io_out_s_21),
    .io_out_s_22(axpy_dp_io_out_s_22),
    .io_out_s_23(axpy_dp_io_out_s_23),
    .io_out_s_24(axpy_dp_io_out_s_24),
    .io_out_s_25(axpy_dp_io_out_s_25),
    .io_out_s_26(axpy_dp_io_out_s_26),
    .io_out_s_27(axpy_dp_io_out_s_27),
    .io_out_s_28(axpy_dp_io_out_s_28),
    .io_out_s_29(axpy_dp_io_out_s_29),
    .io_out_s_30(axpy_dp_io_out_s_30),
    .io_out_s_31(axpy_dp_io_out_s_31),
    .io_out_s_32(axpy_dp_io_out_s_32),
    .io_out_s_33(axpy_dp_io_out_s_33),
    .io_out_s_34(axpy_dp_io_out_s_34),
    .io_out_s_35(axpy_dp_io_out_s_35),
    .io_out_s_36(axpy_dp_io_out_s_36),
    .io_out_s_37(axpy_dp_io_out_s_37),
    .io_out_s_38(axpy_dp_io_out_s_38),
    .io_out_s_39(axpy_dp_io_out_s_39),
    .io_out_s_40(axpy_dp_io_out_s_40),
    .io_out_s_41(axpy_dp_io_out_s_41),
    .io_out_s_42(axpy_dp_io_out_s_42),
    .io_out_s_43(axpy_dp_io_out_s_43),
    .io_out_s_44(axpy_dp_io_out_s_44),
    .io_out_s_45(axpy_dp_io_out_s_45),
    .io_out_s_46(axpy_dp_io_out_s_46),
    .io_out_s_47(axpy_dp_io_out_s_47),
    .io_out_s_48(axpy_dp_io_out_s_48),
    .io_out_s_49(axpy_dp_io_out_s_49),
    .io_out_s_50(axpy_dp_io_out_s_50),
    .io_out_s_51(axpy_dp_io_out_s_51),
    .io_out_s_52(axpy_dp_io_out_s_52),
    .io_out_s_53(axpy_dp_io_out_s_53),
    .io_out_s_54(axpy_dp_io_out_s_54),
    .io_out_s_55(axpy_dp_io_out_s_55),
    .io_out_s_56(axpy_dp_io_out_s_56),
    .io_out_s_57(axpy_dp_io_out_s_57),
    .io_out_s_58(axpy_dp_io_out_s_58),
    .io_out_s_59(axpy_dp_io_out_s_59),
    .io_out_s_60(axpy_dp_io_out_s_60),
    .io_out_s_61(axpy_dp_io_out_s_61),
    .io_out_s_62(axpy_dp_io_out_s_62),
    .io_out_s_63(axpy_dp_io_out_s_63),
    .io_out_s_64(axpy_dp_io_out_s_64),
    .io_out_s_65(axpy_dp_io_out_s_65),
    .io_out_s_66(axpy_dp_io_out_s_66),
    .io_out_s_67(axpy_dp_io_out_s_67),
    .io_out_s_68(axpy_dp_io_out_s_68),
    .io_out_s_69(axpy_dp_io_out_s_69),
    .io_out_s_70(axpy_dp_io_out_s_70),
    .io_out_s_71(axpy_dp_io_out_s_71),
    .io_out_s_72(axpy_dp_io_out_s_72),
    .io_out_s_73(axpy_dp_io_out_s_73),
    .io_out_s_74(axpy_dp_io_out_s_74),
    .io_out_s_75(axpy_dp_io_out_s_75),
    .io_out_s_76(axpy_dp_io_out_s_76),
    .io_out_s_77(axpy_dp_io_out_s_77),
    .io_out_s_78(axpy_dp_io_out_s_78),
    .io_out_s_79(axpy_dp_io_out_s_79),
    .io_out_s_80(axpy_dp_io_out_s_80),
    .io_out_s_81(axpy_dp_io_out_s_81),
    .io_out_s_82(axpy_dp_io_out_s_82),
    .io_out_s_83(axpy_dp_io_out_s_83),
    .io_out_s_84(axpy_dp_io_out_s_84),
    .io_out_s_85(axpy_dp_io_out_s_85),
    .io_out_s_86(axpy_dp_io_out_s_86),
    .io_out_s_87(axpy_dp_io_out_s_87),
    .io_out_s_88(axpy_dp_io_out_s_88),
    .io_out_s_89(axpy_dp_io_out_s_89),
    .io_out_s_90(axpy_dp_io_out_s_90),
    .io_out_s_91(axpy_dp_io_out_s_91),
    .io_out_s_92(axpy_dp_io_out_s_92),
    .io_out_s_93(axpy_dp_io_out_s_93),
    .io_out_s_94(axpy_dp_io_out_s_94),
    .io_out_s_95(axpy_dp_io_out_s_95),
    .io_out_s_96(axpy_dp_io_out_s_96),
    .io_out_s_97(axpy_dp_io_out_s_97),
    .io_out_s_98(axpy_dp_io_out_s_98),
    .io_out_s_99(axpy_dp_io_out_s_99),
    .io_out_s_100(axpy_dp_io_out_s_100),
    .io_out_s_101(axpy_dp_io_out_s_101),
    .io_out_s_102(axpy_dp_io_out_s_102),
    .io_out_s_103(axpy_dp_io_out_s_103),
    .io_out_s_104(axpy_dp_io_out_s_104),
    .io_out_s_105(axpy_dp_io_out_s_105),
    .io_out_s_106(axpy_dp_io_out_s_106),
    .io_out_s_107(axpy_dp_io_out_s_107),
    .io_out_s_108(axpy_dp_io_out_s_108),
    .io_out_s_109(axpy_dp_io_out_s_109),
    .io_out_s_110(axpy_dp_io_out_s_110),
    .io_out_s_111(axpy_dp_io_out_s_111),
    .io_out_s_112(axpy_dp_io_out_s_112),
    .io_out_s_113(axpy_dp_io_out_s_113),
    .io_out_s_114(axpy_dp_io_out_s_114),
    .io_out_s_115(axpy_dp_io_out_s_115),
    .io_out_s_116(axpy_dp_io_out_s_116),
    .io_out_s_117(axpy_dp_io_out_s_117),
    .io_out_s_118(axpy_dp_io_out_s_118),
    .io_out_s_119(axpy_dp_io_out_s_119),
    .io_out_s_120(axpy_dp_io_out_s_120),
    .io_out_s_121(axpy_dp_io_out_s_121),
    .io_out_s_122(axpy_dp_io_out_s_122),
    .io_out_s_123(axpy_dp_io_out_s_123),
    .io_out_s_124(axpy_dp_io_out_s_124),
    .io_out_s_125(axpy_dp_io_out_s_125),
    .io_out_s_126(axpy_dp_io_out_s_126),
    .io_out_s_127(axpy_dp_io_out_s_127)
  );
  assign io_hh_dout = {io_hh_dout_hi,io_hh_dout_lo}; // @[hh_datapath_chisel.scala 286:28]
  assign FP_DDOT_dp_clock = io_clk;
  assign FP_DDOT_dp_reset = io_rst;
  assign FP_DDOT_dp_io_in_a_0 = ddot_din_a[4095:4064]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_1 = ddot_din_a[4063:4032]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_2 = ddot_din_a[4031:4000]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_3 = ddot_din_a[3999:3968]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_4 = ddot_din_a[3967:3936]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_5 = ddot_din_a[3935:3904]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_6 = ddot_din_a[3903:3872]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_7 = ddot_din_a[3871:3840]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_8 = ddot_din_a[3839:3808]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_9 = ddot_din_a[3807:3776]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_10 = ddot_din_a[3775:3744]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_11 = ddot_din_a[3743:3712]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_12 = ddot_din_a[3711:3680]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_13 = ddot_din_a[3679:3648]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_14 = ddot_din_a[3647:3616]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_15 = ddot_din_a[3615:3584]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_16 = ddot_din_a[3583:3552]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_17 = ddot_din_a[3551:3520]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_18 = ddot_din_a[3519:3488]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_19 = ddot_din_a[3487:3456]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_20 = ddot_din_a[3455:3424]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_21 = ddot_din_a[3423:3392]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_22 = ddot_din_a[3391:3360]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_23 = ddot_din_a[3359:3328]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_24 = ddot_din_a[3327:3296]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_25 = ddot_din_a[3295:3264]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_26 = ddot_din_a[3263:3232]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_27 = ddot_din_a[3231:3200]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_28 = ddot_din_a[3199:3168]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_29 = ddot_din_a[3167:3136]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_30 = ddot_din_a[3135:3104]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_31 = ddot_din_a[3103:3072]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_32 = ddot_din_a[3071:3040]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_33 = ddot_din_a[3039:3008]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_34 = ddot_din_a[3007:2976]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_35 = ddot_din_a[2975:2944]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_36 = ddot_din_a[2943:2912]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_37 = ddot_din_a[2911:2880]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_38 = ddot_din_a[2879:2848]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_39 = ddot_din_a[2847:2816]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_40 = ddot_din_a[2815:2784]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_41 = ddot_din_a[2783:2752]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_42 = ddot_din_a[2751:2720]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_43 = ddot_din_a[2719:2688]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_44 = ddot_din_a[2687:2656]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_45 = ddot_din_a[2655:2624]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_46 = ddot_din_a[2623:2592]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_47 = ddot_din_a[2591:2560]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_48 = ddot_din_a[2559:2528]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_49 = ddot_din_a[2527:2496]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_50 = ddot_din_a[2495:2464]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_51 = ddot_din_a[2463:2432]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_52 = ddot_din_a[2431:2400]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_53 = ddot_din_a[2399:2368]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_54 = ddot_din_a[2367:2336]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_55 = ddot_din_a[2335:2304]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_56 = ddot_din_a[2303:2272]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_57 = ddot_din_a[2271:2240]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_58 = ddot_din_a[2239:2208]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_59 = ddot_din_a[2207:2176]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_60 = ddot_din_a[2175:2144]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_61 = ddot_din_a[2143:2112]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_62 = ddot_din_a[2111:2080]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_63 = ddot_din_a[2079:2048]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_64 = ddot_din_a[2047:2016]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_65 = ddot_din_a[2015:1984]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_66 = ddot_din_a[1983:1952]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_67 = ddot_din_a[1951:1920]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_68 = ddot_din_a[1919:1888]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_69 = ddot_din_a[1887:1856]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_70 = ddot_din_a[1855:1824]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_71 = ddot_din_a[1823:1792]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_72 = ddot_din_a[1791:1760]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_73 = ddot_din_a[1759:1728]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_74 = ddot_din_a[1727:1696]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_75 = ddot_din_a[1695:1664]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_76 = ddot_din_a[1663:1632]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_77 = ddot_din_a[1631:1600]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_78 = ddot_din_a[1599:1568]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_79 = ddot_din_a[1567:1536]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_80 = ddot_din_a[1535:1504]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_81 = ddot_din_a[1503:1472]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_82 = ddot_din_a[1471:1440]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_83 = ddot_din_a[1439:1408]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_84 = ddot_din_a[1407:1376]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_85 = ddot_din_a[1375:1344]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_86 = ddot_din_a[1343:1312]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_87 = ddot_din_a[1311:1280]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_88 = ddot_din_a[1279:1248]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_89 = ddot_din_a[1247:1216]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_90 = ddot_din_a[1215:1184]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_91 = ddot_din_a[1183:1152]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_92 = ddot_din_a[1151:1120]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_93 = ddot_din_a[1119:1088]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_94 = ddot_din_a[1087:1056]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_95 = ddot_din_a[1055:1024]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_96 = ddot_din_a[1023:992]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_97 = ddot_din_a[991:960]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_98 = ddot_din_a[959:928]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_99 = ddot_din_a[927:896]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_100 = ddot_din_a[895:864]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_101 = ddot_din_a[863:832]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_102 = ddot_din_a[831:800]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_103 = ddot_din_a[799:768]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_104 = ddot_din_a[767:736]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_105 = ddot_din_a[735:704]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_106 = ddot_din_a[703:672]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_107 = ddot_din_a[671:640]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_108 = ddot_din_a[639:608]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_109 = ddot_din_a[607:576]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_110 = ddot_din_a[575:544]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_111 = ddot_din_a[543:512]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_112 = ddot_din_a[511:480]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_113 = ddot_din_a[479:448]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_114 = ddot_din_a[447:416]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_115 = ddot_din_a[415:384]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_116 = ddot_din_a[383:352]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_117 = ddot_din_a[351:320]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_118 = ddot_din_a[319:288]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_119 = ddot_din_a[287:256]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_120 = ddot_din_a[255:224]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_121 = ddot_din_a[223:192]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_122 = ddot_din_a[191:160]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_123 = ddot_din_a[159:128]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_124 = ddot_din_a[127:96]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_125 = ddot_din_a[95:64]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_126 = ddot_din_a[63:32]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_a_127 = ddot_din_a[31:0]; // @[hh_datapath_chisel.scala 251:33]
  assign FP_DDOT_dp_io_in_b_0 = ddot_din_b[4095:4064]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_1 = ddot_din_b[4063:4032]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_2 = ddot_din_b[4031:4000]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_3 = ddot_din_b[3999:3968]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_4 = ddot_din_b[3967:3936]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_5 = ddot_din_b[3935:3904]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_6 = ddot_din_b[3903:3872]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_7 = ddot_din_b[3871:3840]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_8 = ddot_din_b[3839:3808]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_9 = ddot_din_b[3807:3776]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_10 = ddot_din_b[3775:3744]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_11 = ddot_din_b[3743:3712]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_12 = ddot_din_b[3711:3680]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_13 = ddot_din_b[3679:3648]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_14 = ddot_din_b[3647:3616]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_15 = ddot_din_b[3615:3584]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_16 = ddot_din_b[3583:3552]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_17 = ddot_din_b[3551:3520]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_18 = ddot_din_b[3519:3488]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_19 = ddot_din_b[3487:3456]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_20 = ddot_din_b[3455:3424]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_21 = ddot_din_b[3423:3392]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_22 = ddot_din_b[3391:3360]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_23 = ddot_din_b[3359:3328]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_24 = ddot_din_b[3327:3296]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_25 = ddot_din_b[3295:3264]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_26 = ddot_din_b[3263:3232]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_27 = ddot_din_b[3231:3200]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_28 = ddot_din_b[3199:3168]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_29 = ddot_din_b[3167:3136]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_30 = ddot_din_b[3135:3104]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_31 = ddot_din_b[3103:3072]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_32 = ddot_din_b[3071:3040]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_33 = ddot_din_b[3039:3008]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_34 = ddot_din_b[3007:2976]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_35 = ddot_din_b[2975:2944]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_36 = ddot_din_b[2943:2912]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_37 = ddot_din_b[2911:2880]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_38 = ddot_din_b[2879:2848]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_39 = ddot_din_b[2847:2816]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_40 = ddot_din_b[2815:2784]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_41 = ddot_din_b[2783:2752]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_42 = ddot_din_b[2751:2720]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_43 = ddot_din_b[2719:2688]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_44 = ddot_din_b[2687:2656]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_45 = ddot_din_b[2655:2624]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_46 = ddot_din_b[2623:2592]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_47 = ddot_din_b[2591:2560]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_48 = ddot_din_b[2559:2528]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_49 = ddot_din_b[2527:2496]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_50 = ddot_din_b[2495:2464]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_51 = ddot_din_b[2463:2432]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_52 = ddot_din_b[2431:2400]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_53 = ddot_din_b[2399:2368]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_54 = ddot_din_b[2367:2336]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_55 = ddot_din_b[2335:2304]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_56 = ddot_din_b[2303:2272]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_57 = ddot_din_b[2271:2240]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_58 = ddot_din_b[2239:2208]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_59 = ddot_din_b[2207:2176]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_60 = ddot_din_b[2175:2144]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_61 = ddot_din_b[2143:2112]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_62 = ddot_din_b[2111:2080]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_63 = ddot_din_b[2079:2048]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_64 = ddot_din_b[2047:2016]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_65 = ddot_din_b[2015:1984]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_66 = ddot_din_b[1983:1952]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_67 = ddot_din_b[1951:1920]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_68 = ddot_din_b[1919:1888]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_69 = ddot_din_b[1887:1856]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_70 = ddot_din_b[1855:1824]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_71 = ddot_din_b[1823:1792]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_72 = ddot_din_b[1791:1760]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_73 = ddot_din_b[1759:1728]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_74 = ddot_din_b[1727:1696]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_75 = ddot_din_b[1695:1664]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_76 = ddot_din_b[1663:1632]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_77 = ddot_din_b[1631:1600]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_78 = ddot_din_b[1599:1568]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_79 = ddot_din_b[1567:1536]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_80 = ddot_din_b[1535:1504]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_81 = ddot_din_b[1503:1472]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_82 = ddot_din_b[1471:1440]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_83 = ddot_din_b[1439:1408]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_84 = ddot_din_b[1407:1376]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_85 = ddot_din_b[1375:1344]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_86 = ddot_din_b[1343:1312]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_87 = ddot_din_b[1311:1280]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_88 = ddot_din_b[1279:1248]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_89 = ddot_din_b[1247:1216]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_90 = ddot_din_b[1215:1184]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_91 = ddot_din_b[1183:1152]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_92 = ddot_din_b[1151:1120]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_93 = ddot_din_b[1119:1088]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_94 = ddot_din_b[1087:1056]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_95 = ddot_din_b[1055:1024]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_96 = ddot_din_b[1023:992]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_97 = ddot_din_b[991:960]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_98 = ddot_din_b[959:928]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_99 = ddot_din_b[927:896]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_100 = ddot_din_b[895:864]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_101 = ddot_din_b[863:832]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_102 = ddot_din_b[831:800]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_103 = ddot_din_b[799:768]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_104 = ddot_din_b[767:736]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_105 = ddot_din_b[735:704]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_106 = ddot_din_b[703:672]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_107 = ddot_din_b[671:640]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_108 = ddot_din_b[639:608]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_109 = ddot_din_b[607:576]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_110 = ddot_din_b[575:544]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_111 = ddot_din_b[543:512]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_112 = ddot_din_b[511:480]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_113 = ddot_din_b[479:448]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_114 = ddot_din_b[447:416]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_115 = ddot_din_b[415:384]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_116 = ddot_din_b[383:352]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_117 = ddot_din_b[351:320]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_118 = ddot_din_b[319:288]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_119 = ddot_din_b[287:256]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_120 = ddot_din_b[255:224]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_121 = ddot_din_b[223:192]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_122 = ddot_din_b[191:160]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_123 = ddot_din_b[159:128]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_124 = ddot_din_b[127:96]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_125 = ddot_din_b[95:64]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_126 = ddot_din_b[63:32]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_DDOT_dp_io_in_b_127 = ddot_din_b[31:0]; // @[hh_datapath_chisel.scala 252:33]
  assign FP_square_root_newfpu_clock = io_clk;
  assign FP_square_root_newfpu_reset = io_rst;
  assign FP_square_root_newfpu_io_in_a = io_d1_vld ? ddot_dout : d1_reg; // @[hh_datapath_chisel.scala 171:20 172:10 174:10]
  assign hqr5_clock = io_clk;
  assign hqr5_reset = io_rst;
  assign hqr5_io_in_a = io_d1_rdy ? x1_update : x1_reg; // @[hh_datapath_chisel.scala 183:20 184:10 186:10]
  assign hqr5_io_in_b = io_d2_vld ? d2_update : d2_reg; // @[hh_datapath_chisel.scala 189:20 190:10 192:10]
  assign hqr7_clock = io_clk;
  assign hqr7_reset = io_rst;
  assign hqr7_io_in_a = io_d3_vld ? ddot_dout : d3_reg; // @[hh_datapath_chisel.scala 177:20 178:10 180:10]
  assign FP_multiplier_10ccs_clock = io_clk;
  assign FP_multiplier_10ccs_reset = io_rst;
  assign FP_multiplier_10ccs_io_in_a = io_d5_rdy ? d4_update : d4_reg; // @[hh_datapath_chisel.scala 207:20 208:10 210:10]
  assign FP_multiplier_10ccs_io_in_b = io_tk_vld ? tk_update : tk_reg; // @[hh_datapath_chisel.scala 201:20 202:10 204:10]
  assign axpy_dp_clock = io_clk;
  assign axpy_dp_reset = io_rst;
  assign axpy_dp_io_in_a = io_d5_vld ? d5_update : d5_reg; // @[hh_datapath_chisel.scala 213:20 214:10 216:10]
  assign axpy_dp_io_in_b_0 = vk[4095:4064]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_1 = vk[4063:4032]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_2 = vk[4031:4000]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_3 = vk[3999:3968]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_4 = vk[3967:3936]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_5 = vk[3935:3904]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_6 = vk[3903:3872]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_7 = vk[3871:3840]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_8 = vk[3839:3808]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_9 = vk[3807:3776]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_10 = vk[3775:3744]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_11 = vk[3743:3712]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_12 = vk[3711:3680]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_13 = vk[3679:3648]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_14 = vk[3647:3616]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_15 = vk[3615:3584]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_16 = vk[3583:3552]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_17 = vk[3551:3520]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_18 = vk[3519:3488]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_19 = vk[3487:3456]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_20 = vk[3455:3424]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_21 = vk[3423:3392]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_22 = vk[3391:3360]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_23 = vk[3359:3328]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_24 = vk[3327:3296]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_25 = vk[3295:3264]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_26 = vk[3263:3232]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_27 = vk[3231:3200]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_28 = vk[3199:3168]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_29 = vk[3167:3136]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_30 = vk[3135:3104]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_31 = vk[3103:3072]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_32 = vk[3071:3040]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_33 = vk[3039:3008]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_34 = vk[3007:2976]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_35 = vk[2975:2944]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_36 = vk[2943:2912]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_37 = vk[2911:2880]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_38 = vk[2879:2848]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_39 = vk[2847:2816]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_40 = vk[2815:2784]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_41 = vk[2783:2752]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_42 = vk[2751:2720]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_43 = vk[2719:2688]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_44 = vk[2687:2656]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_45 = vk[2655:2624]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_46 = vk[2623:2592]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_47 = vk[2591:2560]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_48 = vk[2559:2528]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_49 = vk[2527:2496]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_50 = vk[2495:2464]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_51 = vk[2463:2432]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_52 = vk[2431:2400]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_53 = vk[2399:2368]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_54 = vk[2367:2336]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_55 = vk[2335:2304]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_56 = vk[2303:2272]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_57 = vk[2271:2240]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_58 = vk[2239:2208]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_59 = vk[2207:2176]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_60 = vk[2175:2144]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_61 = vk[2143:2112]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_62 = vk[2111:2080]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_63 = vk[2079:2048]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_64 = vk[2047:2016]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_65 = vk[2015:1984]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_66 = vk[1983:1952]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_67 = vk[1951:1920]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_68 = vk[1919:1888]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_69 = vk[1887:1856]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_70 = vk[1855:1824]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_71 = vk[1823:1792]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_72 = vk[1791:1760]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_73 = vk[1759:1728]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_74 = vk[1727:1696]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_75 = vk[1695:1664]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_76 = vk[1663:1632]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_77 = vk[1631:1600]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_78 = vk[1599:1568]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_79 = vk[1567:1536]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_80 = vk[1535:1504]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_81 = vk[1503:1472]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_82 = vk[1471:1440]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_83 = vk[1439:1408]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_84 = vk[1407:1376]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_85 = vk[1375:1344]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_86 = vk[1343:1312]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_87 = vk[1311:1280]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_88 = vk[1279:1248]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_89 = vk[1247:1216]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_90 = vk[1215:1184]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_91 = vk[1183:1152]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_92 = vk[1151:1120]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_93 = vk[1119:1088]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_94 = vk[1087:1056]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_95 = vk[1055:1024]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_96 = vk[1023:992]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_97 = vk[991:960]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_98 = vk[959:928]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_99 = vk[927:896]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_100 = vk[895:864]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_101 = vk[863:832]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_102 = vk[831:800]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_103 = vk[799:768]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_104 = vk[767:736]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_105 = vk[735:704]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_106 = vk[703:672]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_107 = vk[671:640]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_108 = vk[639:608]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_109 = vk[607:576]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_110 = vk[575:544]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_111 = vk[543:512]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_112 = vk[511:480]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_113 = vk[479:448]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_114 = vk[447:416]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_115 = vk[415:384]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_116 = vk[383:352]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_117 = vk[351:320]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_118 = vk[319:288]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_119 = vk[287:256]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_120 = vk[255:224]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_121 = vk[223:192]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_122 = vk[191:160]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_123 = vk[159:128]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_124 = vk[127:96]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_125 = vk[95:64]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_126 = vk[63:32]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_127 = vk[31:0]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_c_0 = yj0[4095:4064]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_1 = yj0[4063:4032]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_2 = yj0[4031:4000]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_3 = yj0[3999:3968]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_4 = yj0[3967:3936]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_5 = yj0[3935:3904]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_6 = yj0[3903:3872]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_7 = yj0[3871:3840]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_8 = yj0[3839:3808]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_9 = yj0[3807:3776]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_10 = yj0[3775:3744]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_11 = yj0[3743:3712]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_12 = yj0[3711:3680]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_13 = yj0[3679:3648]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_14 = yj0[3647:3616]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_15 = yj0[3615:3584]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_16 = yj0[3583:3552]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_17 = yj0[3551:3520]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_18 = yj0[3519:3488]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_19 = yj0[3487:3456]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_20 = yj0[3455:3424]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_21 = yj0[3423:3392]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_22 = yj0[3391:3360]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_23 = yj0[3359:3328]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_24 = yj0[3327:3296]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_25 = yj0[3295:3264]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_26 = yj0[3263:3232]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_27 = yj0[3231:3200]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_28 = yj0[3199:3168]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_29 = yj0[3167:3136]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_30 = yj0[3135:3104]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_31 = yj0[3103:3072]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_32 = yj0[3071:3040]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_33 = yj0[3039:3008]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_34 = yj0[3007:2976]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_35 = yj0[2975:2944]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_36 = yj0[2943:2912]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_37 = yj0[2911:2880]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_38 = yj0[2879:2848]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_39 = yj0[2847:2816]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_40 = yj0[2815:2784]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_41 = yj0[2783:2752]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_42 = yj0[2751:2720]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_43 = yj0[2719:2688]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_44 = yj0[2687:2656]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_45 = yj0[2655:2624]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_46 = yj0[2623:2592]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_47 = yj0[2591:2560]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_48 = yj0[2559:2528]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_49 = yj0[2527:2496]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_50 = yj0[2495:2464]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_51 = yj0[2463:2432]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_52 = yj0[2431:2400]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_53 = yj0[2399:2368]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_54 = yj0[2367:2336]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_55 = yj0[2335:2304]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_56 = yj0[2303:2272]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_57 = yj0[2271:2240]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_58 = yj0[2239:2208]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_59 = yj0[2207:2176]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_60 = yj0[2175:2144]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_61 = yj0[2143:2112]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_62 = yj0[2111:2080]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_63 = yj0[2079:2048]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_64 = yj0[2047:2016]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_65 = yj0[2015:1984]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_66 = yj0[1983:1952]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_67 = yj0[1951:1920]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_68 = yj0[1919:1888]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_69 = yj0[1887:1856]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_70 = yj0[1855:1824]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_71 = yj0[1823:1792]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_72 = yj0[1791:1760]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_73 = yj0[1759:1728]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_74 = yj0[1727:1696]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_75 = yj0[1695:1664]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_76 = yj0[1663:1632]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_77 = yj0[1631:1600]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_78 = yj0[1599:1568]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_79 = yj0[1567:1536]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_80 = yj0[1535:1504]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_81 = yj0[1503:1472]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_82 = yj0[1471:1440]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_83 = yj0[1439:1408]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_84 = yj0[1407:1376]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_85 = yj0[1375:1344]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_86 = yj0[1343:1312]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_87 = yj0[1311:1280]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_88 = yj0[1279:1248]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_89 = yj0[1247:1216]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_90 = yj0[1215:1184]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_91 = yj0[1183:1152]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_92 = yj0[1151:1120]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_93 = yj0[1119:1088]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_94 = yj0[1087:1056]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_95 = yj0[1055:1024]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_96 = yj0[1023:992]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_97 = yj0[991:960]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_98 = yj0[959:928]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_99 = yj0[927:896]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_100 = yj0[895:864]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_101 = yj0[863:832]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_102 = yj0[831:800]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_103 = yj0[799:768]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_104 = yj0[767:736]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_105 = yj0[735:704]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_106 = yj0[703:672]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_107 = yj0[671:640]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_108 = yj0[639:608]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_109 = yj0[607:576]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_110 = yj0[575:544]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_111 = yj0[543:512]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_112 = yj0[511:480]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_113 = yj0[479:448]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_114 = yj0[447:416]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_115 = yj0[415:384]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_116 = yj0[383:352]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_117 = yj0[351:320]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_118 = yj0[319:288]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_119 = yj0[287:256]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_120 = yj0[255:224]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_121 = yj0[223:192]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_122 = yj0[191:160]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_123 = yj0[159:128]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_124 = yj0[127:96]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_125 = yj0[95:64]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_126 = yj0[63:32]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_127 = yj0[31:0]; // @[hh_datapath_chisel.scala 280:26]
  always @(posedge io_clk) begin
    if (io_rst) begin // @[hh_datapath_chisel.scala 59:17]
      yj0 <= 4096'h0; // @[hh_datapath_chisel.scala 64:11]
    end else if (io_yj_sft) begin // @[hh_datapath_chisel.scala 65:26]
      yj0 <= yj_reg_4[4095:0]; // @[hh_datapath_chisel.scala 70:11]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 59:17]
      yj_reg_1 <= 243712'h0; // @[hh_datapath_chisel.scala 60:16]
    end else if (io_yj_sft) begin // @[hh_datapath_chisel.scala 65:26]
      yj_reg_1 <= _yj_reg_1_T[247807:4096]; // @[hh_datapath_chisel.scala 69:16]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 59:17]
      yj_reg_2 <= 243712'h0; // @[hh_datapath_chisel.scala 61:16]
    end else if (io_yj_sft) begin // @[hh_datapath_chisel.scala 65:26]
      yj_reg_2 <= _yj_reg_2_T_1[247807:4096]; // @[hh_datapath_chisel.scala 68:16]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 59:17]
      yj_reg_3 <= 243712'h0; // @[hh_datapath_chisel.scala 62:16]
    end else if (io_yj_sft) begin // @[hh_datapath_chisel.scala 65:26]
      yj_reg_3 <= _yj_reg_3_T_1[247807:4096]; // @[hh_datapath_chisel.scala 67:16]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 59:17]
      yj_reg_4 <= 243712'h0; // @[hh_datapath_chisel.scala 63:16]
    end else if (io_yj_sft) begin // @[hh_datapath_chisel.scala 65:26]
      yj_reg_4 <= _yj_reg_4_T_1[247807:4096]; // @[hh_datapath_chisel.scala 66:16]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      ddot_din_a_reg <= 4096'h0; // @[hh_datapath_chisel.scala 110:22]
    end else if (io_d1_rdy) begin // @[hh_datapath_chisel.scala 135:20]
      ddot_din_a_reg <= io_hh_din; // @[hh_datapath_chisel.scala 136:18]
    end else if (io_d3_rdy) begin // @[hh_datapath_chisel.scala 137:26]
      if (io_vk1_vld) begin // @[hh_datapath_chisel.scala 155:21]
        ddot_din_a_reg <= vk_update; // @[hh_datapath_chisel.scala 156:10]
      end else begin
        ddot_din_a_reg <= vk_reg; // @[hh_datapath_chisel.scala 158:10]
      end
    end else if (io_d4_rdy) begin // @[hh_datapath_chisel.scala 139:26]
      ddot_din_a_reg <= io_hh_din; // @[hh_datapath_chisel.scala 140:18]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      ddot_din_b_reg <= 4096'h0; // @[hh_datapath_chisel.scala 111:22]
    end else if (io_d1_rdy) begin // @[hh_datapath_chisel.scala 145:20]
      ddot_din_b_reg <= io_hh_din; // @[hh_datapath_chisel.scala 146:18]
    end else if (io_d3_rdy) begin // @[hh_datapath_chisel.scala 147:26]
      ddot_din_b_reg <= vk; // @[hh_datapath_chisel.scala 148:18]
    end else if (io_d4_rdy) begin // @[hh_datapath_chisel.scala 149:26]
      ddot_din_b_reg <= vk; // @[hh_datapath_chisel.scala 150:18]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      vk_reg <= 4096'h0; // @[hh_datapath_chisel.scala 112:14]
    end else if (io_vk1_vld) begin // @[hh_datapath_chisel.scala 155:21]
      vk_reg <= vk_update; // @[hh_datapath_chisel.scala 156:10]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      d1_reg <= 32'h0; // @[hh_datapath_chisel.scala 113:14]
    end else if (io_d1_vld) begin // @[hh_datapath_chisel.scala 171:20]
      d1_reg <= ddot_dout; // @[hh_datapath_chisel.scala 172:10]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      d3_reg <= 32'h0; // @[hh_datapath_chisel.scala 114:14]
    end else if (io_d3_vld) begin // @[hh_datapath_chisel.scala 177:20]
      d3_reg <= ddot_dout; // @[hh_datapath_chisel.scala 178:10]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 162:17]
      d4_update <= 32'h0; // @[hh_datapath_chisel.scala 163:17]
    end else if (io_d4_sft) begin // @[hh_datapath_chisel.scala 165:26]
      d4_update <= d4_update_reg[31:0]; // @[hh_datapath_chisel.scala 168:17]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      x1_reg <= 32'h0; // @[hh_datapath_chisel.scala 115:14]
    end else if (io_d1_rdy) begin // @[hh_datapath_chisel.scala 183:20]
      if (io_rst) begin // @[hh_datapath_chisel.scala 223:17]
        x1_reg <= 32'h0; // @[hh_datapath_chisel.scala 224:17]
      end else if (io_d1_rdy) begin // @[hh_datapath_chisel.scala 225:26]
        x1_reg <= _GEN_167; // @[hh_datapath_chisel.scala 226:17]
      end else begin
        x1_reg <= 32'h0; // @[hh_datapath_chisel.scala 228:17]
      end
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      d2_reg <= 32'h0; // @[hh_datapath_chisel.scala 116:14]
    end else if (io_d2_vld) begin // @[hh_datapath_chisel.scala 189:20]
      d2_reg <= d2_update; // @[hh_datapath_chisel.scala 190:10]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      vk1_reg <= 32'h0; // @[hh_datapath_chisel.scala 117:15]
    end else if (io_vk1_vld) begin // @[hh_datapath_chisel.scala 195:21]
      vk1_reg <= vk1_update; // @[hh_datapath_chisel.scala 196:11]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      tk_reg <= 32'h0; // @[hh_datapath_chisel.scala 118:14]
    end else if (io_tk_vld) begin // @[hh_datapath_chisel.scala 201:20]
      tk_reg <= tk_update; // @[hh_datapath_chisel.scala 202:10]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      d4_reg <= 32'h0; // @[hh_datapath_chisel.scala 119:14]
    end else if (io_d5_rdy) begin // @[hh_datapath_chisel.scala 207:20]
      d4_reg <= d4_update; // @[hh_datapath_chisel.scala 208:10]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      d5_reg <= 32'h0; // @[hh_datapath_chisel.scala 120:14]
    end else if (io_d5_vld) begin // @[hh_datapath_chisel.scala 213:20]
      d5_reg <= d5_update; // @[hh_datapath_chisel.scala 214:10]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 162:17]
      d4_update_reg <= 4064'h0; // @[hh_datapath_chisel.scala 164:21]
    end else if (io_d4_sft) begin // @[hh_datapath_chisel.scala 165:26]
      d4_update_reg <= _d4_update_reg_T[4095:32]; // @[hh_datapath_chisel.scala 167:21]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {128{`RANDOM}};
  yj0 = _RAND_0[4095:0];
  _RAND_1 = {7616{`RANDOM}};
  yj_reg_1 = _RAND_1[243711:0];
  _RAND_2 = {7616{`RANDOM}};
  yj_reg_2 = _RAND_2[243711:0];
  _RAND_3 = {7616{`RANDOM}};
  yj_reg_3 = _RAND_3[243711:0];
  _RAND_4 = {7616{`RANDOM}};
  yj_reg_4 = _RAND_4[243711:0];
  _RAND_5 = {128{`RANDOM}};
  ddot_din_a_reg = _RAND_5[4095:0];
  _RAND_6 = {128{`RANDOM}};
  ddot_din_b_reg = _RAND_6[4095:0];
  _RAND_7 = {128{`RANDOM}};
  vk_reg = _RAND_7[4095:0];
  _RAND_8 = {1{`RANDOM}};
  d1_reg = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  d3_reg = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  d4_update = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  x1_reg = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  d2_reg = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  vk1_reg = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  tk_reg = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  d4_reg = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  d5_reg = _RAND_16[31:0];
  _RAND_17 = {127{`RANDOM}};
  d4_update_reg = _RAND_17[4063:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module hh_datapath(
  input           clk,
  input           rst,
  input  [15:0]   hh_cnt,
  input           d1_rdy,
  input           d1_vld,
  input           d2_rdy,
  input           d2_vld,
  input           vk1_rdy,
  input           vk1_vld,
  input           d3_rdy,
  input           d3_vld,
  input           tk_rdy,
  input           tk_vld,
  input           d4_rdy,
  input           d4_vld,
  input           d5_rdy,
  input           d5_vld,
  input           yjp_rdy,
  input           yjp_vld,
  input           yj_sft,
  input           d4_sft,
  input  [4095:0] hh_din,
  output [4095:0] hh_dout
);
  wire  hh_datapath_1_io_clk; // @[hh_datapath_chisel.scala 315:62]
  wire  hh_datapath_1_io_rst; // @[hh_datapath_chisel.scala 315:62]
  wire [15:0] hh_datapath_1_io_hh_cnt; // @[hh_datapath_chisel.scala 315:62]
  wire  hh_datapath_1_io_d1_rdy; // @[hh_datapath_chisel.scala 315:62]
  wire  hh_datapath_1_io_d1_vld; // @[hh_datapath_chisel.scala 315:62]
  wire  hh_datapath_1_io_d2_vld; // @[hh_datapath_chisel.scala 315:62]
  wire  hh_datapath_1_io_vk1_vld; // @[hh_datapath_chisel.scala 315:62]
  wire  hh_datapath_1_io_d3_rdy; // @[hh_datapath_chisel.scala 315:62]
  wire  hh_datapath_1_io_d3_vld; // @[hh_datapath_chisel.scala 315:62]
  wire  hh_datapath_1_io_tk_vld; // @[hh_datapath_chisel.scala 315:62]
  wire  hh_datapath_1_io_d4_rdy; // @[hh_datapath_chisel.scala 315:62]
  wire  hh_datapath_1_io_d5_rdy; // @[hh_datapath_chisel.scala 315:62]
  wire  hh_datapath_1_io_d5_vld; // @[hh_datapath_chisel.scala 315:62]
  wire  hh_datapath_1_io_yj_sft; // @[hh_datapath_chisel.scala 315:62]
  wire  hh_datapath_1_io_d4_sft; // @[hh_datapath_chisel.scala 315:62]
  wire [4095:0] hh_datapath_1_io_hh_din; // @[hh_datapath_chisel.scala 315:62]
  wire [4095:0] hh_datapath_1_io_hh_dout; // @[hh_datapath_chisel.scala 315:62]
  hh_datapath_1 hh_datapath_1 ( // @[hh_datapath_chisel.scala 315:62]
    .io_clk(hh_datapath_1_io_clk),
    .io_rst(hh_datapath_1_io_rst),
    .io_hh_cnt(hh_datapath_1_io_hh_cnt),
    .io_d1_rdy(hh_datapath_1_io_d1_rdy),
    .io_d1_vld(hh_datapath_1_io_d1_vld),
    .io_d2_vld(hh_datapath_1_io_d2_vld),
    .io_vk1_vld(hh_datapath_1_io_vk1_vld),
    .io_d3_rdy(hh_datapath_1_io_d3_rdy),
    .io_d3_vld(hh_datapath_1_io_d3_vld),
    .io_tk_vld(hh_datapath_1_io_tk_vld),
    .io_d4_rdy(hh_datapath_1_io_d4_rdy),
    .io_d5_rdy(hh_datapath_1_io_d5_rdy),
    .io_d5_vld(hh_datapath_1_io_d5_vld),
    .io_yj_sft(hh_datapath_1_io_yj_sft),
    .io_d4_sft(hh_datapath_1_io_d4_sft),
    .io_hh_din(hh_datapath_1_io_hh_din),
    .io_hh_dout(hh_datapath_1_io_hh_dout)
  );
  assign hh_dout = hh_datapath_1_io_hh_dout; // @[hh_datapath_chisel.scala 338:17]
  assign hh_datapath_1_io_clk = clk; // @[hh_datapath_chisel.scala 316:30]
  assign hh_datapath_1_io_rst = rst; // @[hh_datapath_chisel.scala 317:30]
  assign hh_datapath_1_io_hh_cnt = hh_cnt; // @[hh_datapath_chisel.scala 318:33]
  assign hh_datapath_1_io_d1_rdy = d1_rdy; // @[hh_datapath_chisel.scala 319:33]
  assign hh_datapath_1_io_d1_vld = d1_vld; // @[hh_datapath_chisel.scala 320:33]
  assign hh_datapath_1_io_d2_vld = d2_vld; // @[hh_datapath_chisel.scala 322:33]
  assign hh_datapath_1_io_vk1_vld = vk1_vld; // @[hh_datapath_chisel.scala 324:34]
  assign hh_datapath_1_io_d3_rdy = d3_rdy; // @[hh_datapath_chisel.scala 325:33]
  assign hh_datapath_1_io_d3_vld = d3_vld; // @[hh_datapath_chisel.scala 326:33]
  assign hh_datapath_1_io_tk_vld = tk_vld; // @[hh_datapath_chisel.scala 328:33]
  assign hh_datapath_1_io_d4_rdy = d4_rdy; // @[hh_datapath_chisel.scala 329:33]
  assign hh_datapath_1_io_d5_rdy = d5_rdy; // @[hh_datapath_chisel.scala 331:33]
  assign hh_datapath_1_io_d5_vld = d5_vld; // @[hh_datapath_chisel.scala 332:33]
  assign hh_datapath_1_io_yj_sft = yj_sft; // @[hh_datapath_chisel.scala 335:33]
  assign hh_datapath_1_io_d4_sft = d4_sft; // @[hh_datapath_chisel.scala 336:33]
  assign hh_datapath_1_io_hh_din = hh_din; // @[hh_datapath_chisel.scala 337:33]
endmodule

